
module openMSP430(aclk, aclk_en, dbg_freeze, dbg_i2c_sda_out, dbg_uart_txd, dco_enable, dco_wkup, dmem_addr_0_, dmem_addr_1_, dmem_addr_2_, dmem_addr_3_, dmem_addr_4_, dmem_addr_5_, dmem_addr_6_, dmem_addr_7_, dmem_addr_8_, dmem_addr_9_, dmem_addr_10_, dmem_addr_11_, dmem_addr_12_, dmem_cen
, dmem_din_0_, dmem_din_1_, dmem_din_2_, dmem_din_3_, dmem_din_4_, dmem_din_5_, dmem_din_6_, dmem_din_7_, dmem_din_8_, dmem_din_9_, dmem_din_10_, dmem_din_11_, dmem_din_12_, dmem_din_13_, dmem_din_14_, dmem_din_15_, dmem_wen_0_, dmem_wen_1_, irq_acc_0_, irq_acc_1_, irq_acc_2_
, irq_acc_3_, irq_acc_4_, irq_acc_5_, irq_acc_6_, irq_acc_7_, irq_acc_8_, irq_acc_9_, irq_acc_10_, irq_acc_11_, irq_acc_12_, irq_acc_13_, lfxt_enable, lfxt_wkup, mclk, dma_dout_0_, dma_dout_1_, dma_dout_2_, dma_dout_3_, dma_dout_4_, dma_dout_5_, dma_dout_6_
, dma_dout_7_, dma_dout_8_, dma_dout_9_, dma_dout_10_, dma_dout_11_, dma_dout_12_, dma_dout_13_, dma_dout_14_, dma_dout_15_, dma_ready, dma_resp, per_addr_0_, per_addr_1_, per_addr_2_, per_addr_3_, per_addr_4_, per_addr_5_, per_addr_6_, per_addr_7_, per_addr_8_, per_addr_9_
, per_addr_10_, per_addr_11_, per_addr_12_, per_addr_13_, per_din_0_, per_din_1_, per_din_2_, per_din_3_, per_din_4_, per_din_5_, per_din_6_, per_din_7_, per_din_8_, per_din_9_, per_din_10_, per_din_11_, per_din_12_, per_din_13_, per_din_14_, per_din_15_, per_en
, per_we_0_, per_we_1_, pmem_addr_0_, pmem_addr_1_, pmem_addr_2_, pmem_addr_3_, pmem_addr_4_, pmem_addr_5_, pmem_addr_6_, pmem_addr_7_, pmem_addr_8_, pmem_addr_9_, pmem_addr_10_, pmem_addr_11_, pmem_addr_12_, pmem_addr_13_, pmem_cen, pmem_din_0_, pmem_din_1_, pmem_din_2_, pmem_din_3_
, pmem_din_4_, pmem_din_5_, pmem_din_6_, pmem_din_7_, pmem_din_8_, pmem_din_9_, pmem_din_10_, pmem_din_11_, pmem_din_12_, pmem_din_13_, pmem_din_14_, pmem_din_15_, pmem_wen_0_, pmem_wen_1_, puc_rst, smclk, smclk_en, cpu_en, dbg_en, dbg_i2c_addr_0_, dbg_i2c_addr_1_
, dbg_i2c_addr_2_, dbg_i2c_addr_3_, dbg_i2c_addr_4_, dbg_i2c_addr_5_, dbg_i2c_addr_6_, dbg_i2c_broadcast_0_, dbg_i2c_broadcast_1_, dbg_i2c_broadcast_2_, dbg_i2c_broadcast_3_, dbg_i2c_broadcast_4_, dbg_i2c_broadcast_5_, dbg_i2c_broadcast_6_, dbg_i2c_scl, dbg_i2c_sda_in, dbg_uart_rxd, dco_clk, dmem_dout_0_, dmem_dout_1_, dmem_dout_2_, dmem_dout_3_, dmem_dout_4_
, dmem_dout_5_, dmem_dout_6_, dmem_dout_7_, dmem_dout_8_, dmem_dout_9_, dmem_dout_10_, dmem_dout_11_, dmem_dout_12_, dmem_dout_13_, dmem_dout_14_, dmem_dout_15_, irq_0_, irq_1_, irq_2_, irq_3_, irq_4_, irq_5_, irq_6_, irq_7_, irq_8_, irq_9_
, irq_10_, irq_11_, irq_12_, irq_13_, lfxt_clk, dma_addr_1_, dma_addr_2_, dma_addr_3_, dma_addr_4_, dma_addr_5_, dma_addr_6_, dma_addr_7_, dma_addr_8_, dma_addr_9_, dma_addr_10_, dma_addr_11_, dma_addr_12_, dma_addr_13_, dma_addr_14_, dma_addr_15_, dma_din_0_
, dma_din_1_, dma_din_2_, dma_din_3_, dma_din_4_, dma_din_5_, dma_din_6_, dma_din_7_, dma_din_8_, dma_din_9_, dma_din_10_, dma_din_11_, dma_din_12_, dma_din_13_, dma_din_14_, dma_din_15_, dma_en, dma_priority, dma_we_0_, dma_we_1_, dma_wkup, nmi
, per_dout_0_, per_dout_1_, per_dout_2_, per_dout_3_, per_dout_4_, per_dout_5_, per_dout_6_, per_dout_7_, per_dout_8_, per_dout_9_, per_dout_10_, per_dout_11_, per_dout_12_, per_dout_13_, per_dout_14_, per_dout_15_, pmem_dout_0_, pmem_dout_1_, pmem_dout_2_, pmem_dout_3_, pmem_dout_4_
, pmem_dout_5_, pmem_dout_6_, pmem_dout_7_, pmem_dout_8_, pmem_dout_9_, pmem_dout_10_, pmem_dout_11_, pmem_dout_12_, pmem_dout_13_, pmem_dout_14_, pmem_dout_15_, reset_n, scan_enable, scan_mode, wkup);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  output aclk;
  wire aclk;
  output aclk_en;
  wire aclk_en;
  wire  clock_module_0.UNUSED_cpuoff ;
  wire  clock_module_0.aclk_div_0_ ;
  wire  clock_module_0.aclk_div_1_ ;
  wire  clock_module_0.aclk_div_2_ ;
  wire  clock_module_0.bcsctl1_4_ ;
  wire  clock_module_0.bcsctl1_5_ ;
  wire  clock_module_0.bcsctl1_rd_12_ ;
  wire  clock_module_0.bcsctl1_rd_13_ ;
  wire  clock_module_0.bcsctl2_1_ ;
  wire  clock_module_0.bcsctl2_2_ ;
  wire  clock_module_0.bcsctl2_3_ ;
  wire  clock_module_0.bcsctl2_rd_1_ ;
  wire  clock_module_0.bcsctl2_rd_2_ ;
  wire  clock_module_0.bcsctl2_rd_3_ ;
  wire  clock_module_0.dbg_cpu_reset ;
  wire  clock_module_0.dbg_rst ;
  wire  clock_module_0.dbg_rst_nxt ;
  wire  clock_module_0.lfxt_clk_dly ;
  wire  clock_module_0.lfxt_clk_s ;
  wire  clock_module_0.oscoff ;
  wire  clock_module_0.por ;
  wire  clock_module_0.por_a ;
  wire  clock_module_0.puc_a ;
  wire  clock_module_0.puc_noscan_n ;
  wire  clock_module_0.scg1 ;
  wire  clock_module_0.smclk_div_0_ ;
  wire  clock_module_0.smclk_div_1_ ;
  wire  clock_module_0.smclk_div_2_ ;
  wire  clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ;
  wire  clock_module_0.sync_cell_puc.data_in ;
  wire  clock_module_0.sync_cell_puc.data_sync_0_ ;
  wire  clock_module_0.sync_reset_por.data_sync_0_ ;
  wire  clock_module_0.wdt_reset ;
  input cpu_en;
  wire cpu_en;
  wire  dbg_0.UNUSED_eu_mab_0_ ;
  wire  dbg_0.UNUSED_eu_mab_10_ ;
  wire  dbg_0.UNUSED_eu_mab_11_ ;
  wire  dbg_0.UNUSED_eu_mab_12_ ;
  wire  dbg_0.UNUSED_eu_mab_13_ ;
  wire  dbg_0.UNUSED_eu_mab_14_ ;
  wire  dbg_0.UNUSED_eu_mab_15_ ;
  wire  dbg_0.UNUSED_eu_mab_1_ ;
  wire  dbg_0.UNUSED_eu_mab_2_ ;
  wire  dbg_0.UNUSED_eu_mab_3_ ;
  wire  dbg_0.UNUSED_eu_mab_4_ ;
  wire  dbg_0.UNUSED_eu_mab_5_ ;
  wire  dbg_0.UNUSED_eu_mab_6_ ;
  wire  dbg_0.UNUSED_eu_mab_7_ ;
  wire  dbg_0.UNUSED_eu_mab_8_ ;
  wire  dbg_0.UNUSED_eu_mab_9_ ;
  wire  dbg_0.UNUSED_eu_mb_en ;
  wire  dbg_0.UNUSED_eu_mb_wr_0_ ;
  wire  dbg_0.UNUSED_eu_mb_wr_1_ ;
  wire  dbg_0.UNUSED_pc_0_ ;
  wire  dbg_0.UNUSED_pc_10_ ;
  wire  dbg_0.UNUSED_pc_11_ ;
  wire  dbg_0.UNUSED_pc_12_ ;
  wire  dbg_0.UNUSED_pc_13_ ;
  wire  dbg_0.UNUSED_pc_14_ ;
  wire  dbg_0.UNUSED_pc_15_ ;
  wire  dbg_0.UNUSED_pc_1_ ;
  wire  dbg_0.UNUSED_pc_2_ ;
  wire  dbg_0.UNUSED_pc_3_ ;
  wire  dbg_0.UNUSED_pc_4_ ;
  wire  dbg_0.UNUSED_pc_5_ ;
  wire  dbg_0.UNUSED_pc_6_ ;
  wire  dbg_0.UNUSED_pc_7_ ;
  wire  dbg_0.UNUSED_pc_8_ ;
  wire  dbg_0.UNUSED_pc_9_ ;
  wire  dbg_0.cpu_ctl_3_ ;
  wire  dbg_0.cpu_ctl_4_ ;
  wire  dbg_0.cpu_ctl_5_ ;
  wire  dbg_0.cpu_stat_2_ ;
  wire  dbg_0.cpu_stat_3_ ;
  wire  dbg_0.cpu_stat_full_0_ ;
  wire  dbg_0.dbg_addr_0_ ;
  wire  dbg_0.dbg_addr_1_ ;
  wire  dbg_0.dbg_addr_2_ ;
  wire  dbg_0.dbg_addr_3_ ;
  wire  dbg_0.dbg_addr_4_ ;
  wire  dbg_0.dbg_addr_5_ ;
  wire  dbg_0.dbg_din_0_ ;
  wire  dbg_0.dbg_din_10_ ;
  wire  dbg_0.dbg_din_11_ ;
  wire  dbg_0.dbg_din_12_ ;
  wire  dbg_0.dbg_din_13_ ;
  wire  dbg_0.dbg_din_14_ ;
  wire  dbg_0.dbg_din_15_ ;
  wire  dbg_0.dbg_din_1_ ;
  wire  dbg_0.dbg_din_2_ ;
  wire  dbg_0.dbg_din_3_ ;
  wire  dbg_0.dbg_din_4_ ;
  wire  dbg_0.dbg_din_5_ ;
  wire  dbg_0.dbg_din_6_ ;
  wire  dbg_0.dbg_din_7_ ;
  wire  dbg_0.dbg_din_8_ ;
  wire  dbg_0.dbg_din_9_ ;
  wire  dbg_0.dbg_dout_0_ ;
  wire  dbg_0.dbg_dout_10_ ;
  wire  dbg_0.dbg_dout_11_ ;
  wire  dbg_0.dbg_dout_12_ ;
  wire  dbg_0.dbg_dout_13_ ;
  wire  dbg_0.dbg_dout_14_ ;
  wire  dbg_0.dbg_dout_15_ ;
  wire  dbg_0.dbg_dout_1_ ;
  wire  dbg_0.dbg_dout_2_ ;
  wire  dbg_0.dbg_dout_3_ ;
  wire  dbg_0.dbg_dout_4_ ;
  wire  dbg_0.dbg_dout_5_ ;
  wire  dbg_0.dbg_dout_6_ ;
  wire  dbg_0.dbg_dout_7_ ;
  wire  dbg_0.dbg_dout_8_ ;
  wire  dbg_0.dbg_dout_9_ ;
  wire  dbg_0.dbg_halt_cmd ;
  wire  dbg_0.dbg_i2c_0.dbg_bw ;
  wire  dbg_0.dbg_i2c_0.dbg_rd ;
  wire  dbg_0.dbg_i2c_0.dbg_state_0_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_1_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_2_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_nxt_0_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_nxt_1_ ;
  wire  dbg_0.dbg_i2c_0.dbg_state_nxt_2_ ;
  wire  dbg_0.dbg_i2c_0.dbg_wr ;
  wire  dbg_0.dbg_i2c_0.i2c_active_seq ;
  wire  dbg_0.dbg_i2c_0.i2c_state_0_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_1_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_2_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_nxt_0_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_nxt_1_ ;
  wire  dbg_0.dbg_i2c_0.i2c_state_nxt_2_ ;
  wire  dbg_0.dbg_i2c_0.mem_burst ;
  wire  dbg_0.dbg_i2c_0.mem_burst_end ;
  wire  dbg_0.dbg_i2c_0.mem_burst_rd ;
  wire  dbg_0.dbg_i2c_0.mem_burst_wr ;
  wire  dbg_0.dbg_i2c_0.mem_bw ;
  wire  dbg_0.dbg_i2c_0.scl ;
  wire  dbg_0.dbg_i2c_0.scl_buf_0_ ;
  wire  dbg_0.dbg_i2c_0.scl_buf_1_ ;
  wire  dbg_0.dbg_i2c_0.scl_dly ;
  wire  dbg_0.dbg_i2c_0.scl_re ;
  wire  dbg_0.dbg_i2c_0.scl_re_dly_0_ ;
  wire  dbg_0.dbg_i2c_0.scl_re_dly_1_ ;
  wire  dbg_0.dbg_i2c_0.scl_sync ;
  wire  dbg_0.dbg_i2c_0.scl_sync_n ;
  wire  dbg_0.dbg_i2c_0.sda_in ;
  wire  dbg_0.dbg_i2c_0.sda_in_buf_0_ ;
  wire  dbg_0.dbg_i2c_0.sda_in_buf_1_ ;
  wire  dbg_0.dbg_i2c_0.sda_in_dly ;
  wire  dbg_0.dbg_i2c_0.sda_in_sync ;
  wire  dbg_0.dbg_i2c_0.sda_in_sync_n ;
  wire  dbg_0.dbg_i2c_0.shift_buf_0_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_1_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_2_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_3_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_4_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_5_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_6_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_7_ ;
  wire  dbg_0.dbg_i2c_0.shift_buf_8_ ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ;
  wire  dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ;
  wire  dbg_0.dbg_mem_addr_0_ ;
  wire  dbg_0.dbg_mem_addr_10_ ;
  wire  dbg_0.dbg_mem_addr_11_ ;
  wire  dbg_0.dbg_mem_addr_12_ ;
  wire  dbg_0.dbg_mem_addr_13_ ;
  wire  dbg_0.dbg_mem_addr_14_ ;
  wire  dbg_0.dbg_mem_addr_15_ ;
  wire  dbg_0.dbg_mem_addr_1_ ;
  wire  dbg_0.dbg_mem_addr_2_ ;
  wire  dbg_0.dbg_mem_addr_3_ ;
  wire  dbg_0.dbg_mem_addr_4_ ;
  wire  dbg_0.dbg_mem_addr_5_ ;
  wire  dbg_0.dbg_mem_addr_6_ ;
  wire  dbg_0.dbg_mem_addr_7_ ;
  wire  dbg_0.dbg_mem_addr_8_ ;
  wire  dbg_0.dbg_mem_addr_9_ ;
  wire  dbg_0.dbg_mem_din_0_ ;
  wire  dbg_0.dbg_mem_din_10_ ;
  wire  dbg_0.dbg_mem_din_11_ ;
  wire  dbg_0.dbg_mem_din_12_ ;
  wire  dbg_0.dbg_mem_din_13_ ;
  wire  dbg_0.dbg_mem_din_14_ ;
  wire  dbg_0.dbg_mem_din_15_ ;
  wire  dbg_0.dbg_mem_din_1_ ;
  wire  dbg_0.dbg_mem_din_2_ ;
  wire  dbg_0.dbg_mem_din_3_ ;
  wire  dbg_0.dbg_mem_din_4_ ;
  wire  dbg_0.dbg_mem_din_5_ ;
  wire  dbg_0.dbg_mem_din_6_ ;
  wire  dbg_0.dbg_mem_din_7_ ;
  wire  dbg_0.dbg_mem_din_8_ ;
  wire  dbg_0.dbg_mem_din_9_ ;
  wire  dbg_0.dbg_mem_en ;
  wire  dbg_0.dbg_mem_rd ;
  wire  dbg_0.dbg_mem_rd_dly ;
  wire  dbg_0.dbg_mem_wr_0_ ;
  wire  dbg_0.dbg_mem_wr_1_ ;
  wire  dbg_0.dbg_rd_rdy ;
  wire  dbg_0.dbg_reg_din_0_ ;
  wire  dbg_0.dbg_reg_din_10_ ;
  wire  dbg_0.dbg_reg_din_11_ ;
  wire  dbg_0.dbg_reg_din_12_ ;
  wire  dbg_0.dbg_reg_din_13_ ;
  wire  dbg_0.dbg_reg_din_14_ ;
  wire  dbg_0.dbg_reg_din_15_ ;
  wire  dbg_0.dbg_reg_din_1_ ;
  wire  dbg_0.dbg_reg_din_2_ ;
  wire  dbg_0.dbg_reg_din_3_ ;
  wire  dbg_0.dbg_reg_din_4_ ;
  wire  dbg_0.dbg_reg_din_5_ ;
  wire  dbg_0.dbg_reg_din_6_ ;
  wire  dbg_0.dbg_reg_din_7_ ;
  wire  dbg_0.dbg_reg_din_8_ ;
  wire  dbg_0.dbg_reg_din_9_ ;
  wire  dbg_0.dbg_reg_wr ;
  wire  dbg_0.decode_noirq ;
  wire  dbg_0.fe_mdb_in_0_ ;
  wire  dbg_0.fe_mdb_in_10_ ;
  wire  dbg_0.fe_mdb_in_11_ ;
  wire  dbg_0.fe_mdb_in_12_ ;
  wire  dbg_0.fe_mdb_in_13_ ;
  wire  dbg_0.fe_mdb_in_14_ ;
  wire  dbg_0.fe_mdb_in_15_ ;
  wire  dbg_0.fe_mdb_in_1_ ;
  wire  dbg_0.fe_mdb_in_2_ ;
  wire  dbg_0.fe_mdb_in_3_ ;
  wire  dbg_0.fe_mdb_in_4_ ;
  wire  dbg_0.fe_mdb_in_5_ ;
  wire  dbg_0.fe_mdb_in_6_ ;
  wire  dbg_0.fe_mdb_in_7_ ;
  wire  dbg_0.fe_mdb_in_8_ ;
  wire  dbg_0.fe_mdb_in_9_ ;
  wire  dbg_0.halt_flag ;
  wire  dbg_0.inc_step_0_ ;
  wire  dbg_0.inc_step_1_ ;
  wire  dbg_0.istep ;
  wire  dbg_0.mem_cnt_0_ ;
  wire  dbg_0.mem_cnt_10_ ;
  wire  dbg_0.mem_cnt_11_ ;
  wire  dbg_0.mem_cnt_12_ ;
  wire  dbg_0.mem_cnt_13_ ;
  wire  dbg_0.mem_cnt_14_ ;
  wire  dbg_0.mem_cnt_15_ ;
  wire  dbg_0.mem_cnt_1_ ;
  wire  dbg_0.mem_cnt_2_ ;
  wire  dbg_0.mem_cnt_3_ ;
  wire  dbg_0.mem_cnt_4_ ;
  wire  dbg_0.mem_cnt_5_ ;
  wire  dbg_0.mem_cnt_6_ ;
  wire  dbg_0.mem_cnt_7_ ;
  wire  dbg_0.mem_cnt_8_ ;
  wire  dbg_0.mem_cnt_9_ ;
  wire  dbg_0.mem_ctl_1_ ;
  wire  dbg_0.mem_ctl_2_ ;
  wire  dbg_0.mem_data_0_ ;
  wire  dbg_0.mem_data_10_ ;
  wire  dbg_0.mem_data_11_ ;
  wire  dbg_0.mem_data_12_ ;
  wire  dbg_0.mem_data_13_ ;
  wire  dbg_0.mem_data_14_ ;
  wire  dbg_0.mem_data_15_ ;
  wire  dbg_0.mem_data_1_ ;
  wire  dbg_0.mem_data_2_ ;
  wire  dbg_0.mem_data_3_ ;
  wire  dbg_0.mem_data_4_ ;
  wire  dbg_0.mem_data_5_ ;
  wire  dbg_0.mem_data_6_ ;
  wire  dbg_0.mem_data_7_ ;
  wire  dbg_0.mem_data_8_ ;
  wire  dbg_0.mem_data_9_ ;
  wire  dbg_0.mem_start ;
  wire  dbg_0.mem_startb ;
  wire  dbg_0.mem_state_0_ ;
  wire  dbg_0.mem_state_1_ ;
  wire  dbg_0.mem_state_nxt_0_ ;
  wire  dbg_0.mem_state_nxt_1_ ;
  input dbg_en;
  wire dbg_en;
  output dbg_freeze;
  wire dbg_freeze;
  input dbg_i2c_addr_0_;
  wire dbg_i2c_addr_0_;
  input dbg_i2c_addr_1_;
  wire dbg_i2c_addr_1_;
  input dbg_i2c_addr_2_;
  wire dbg_i2c_addr_2_;
  input dbg_i2c_addr_3_;
  wire dbg_i2c_addr_3_;
  input dbg_i2c_addr_4_;
  wire dbg_i2c_addr_4_;
  input dbg_i2c_addr_5_;
  wire dbg_i2c_addr_5_;
  input dbg_i2c_addr_6_;
  wire dbg_i2c_addr_6_;
  input dbg_i2c_broadcast_0_;
  wire dbg_i2c_broadcast_0_;
  input dbg_i2c_broadcast_1_;
  wire dbg_i2c_broadcast_1_;
  input dbg_i2c_broadcast_2_;
  wire dbg_i2c_broadcast_2_;
  input dbg_i2c_broadcast_3_;
  wire dbg_i2c_broadcast_3_;
  input dbg_i2c_broadcast_4_;
  wire dbg_i2c_broadcast_4_;
  input dbg_i2c_broadcast_5_;
  wire dbg_i2c_broadcast_5_;
  input dbg_i2c_broadcast_6_;
  wire dbg_i2c_broadcast_6_;
  input dbg_i2c_scl;
  wire dbg_i2c_scl;
  input dbg_i2c_sda_in;
  wire dbg_i2c_sda_in;
  output dbg_i2c_sda_out;
  wire dbg_i2c_sda_out;
  input dbg_uart_rxd;
  wire dbg_uart_rxd;
  output dbg_uart_txd;
  wire dbg_uart_txd;
  input dco_clk;
  wire dco_clk;
  output dco_enable;
  wire dco_enable;
  output dco_wkup;
  wire dco_wkup;
  input dma_addr_10_;
  wire dma_addr_10_;
  input dma_addr_11_;
  wire dma_addr_11_;
  input dma_addr_12_;
  wire dma_addr_12_;
  input dma_addr_13_;
  wire dma_addr_13_;
  input dma_addr_14_;
  wire dma_addr_14_;
  input dma_addr_15_;
  wire dma_addr_15_;
  input dma_addr_1_;
  wire dma_addr_1_;
  input dma_addr_2_;
  wire dma_addr_2_;
  input dma_addr_3_;
  wire dma_addr_3_;
  input dma_addr_4_;
  wire dma_addr_4_;
  input dma_addr_5_;
  wire dma_addr_5_;
  input dma_addr_6_;
  wire dma_addr_6_;
  input dma_addr_7_;
  wire dma_addr_7_;
  input dma_addr_8_;
  wire dma_addr_8_;
  input dma_addr_9_;
  wire dma_addr_9_;
  input dma_din_0_;
  wire dma_din_0_;
  input dma_din_10_;
  wire dma_din_10_;
  input dma_din_11_;
  wire dma_din_11_;
  input dma_din_12_;
  wire dma_din_12_;
  input dma_din_13_;
  wire dma_din_13_;
  input dma_din_14_;
  wire dma_din_14_;
  input dma_din_15_;
  wire dma_din_15_;
  input dma_din_1_;
  wire dma_din_1_;
  input dma_din_2_;
  wire dma_din_2_;
  input dma_din_3_;
  wire dma_din_3_;
  input dma_din_4_;
  wire dma_din_4_;
  input dma_din_5_;
  wire dma_din_5_;
  input dma_din_6_;
  wire dma_din_6_;
  input dma_din_7_;
  wire dma_din_7_;
  input dma_din_8_;
  wire dma_din_8_;
  input dma_din_9_;
  wire dma_din_9_;
  output dma_dout_0_;
  wire dma_dout_0_;
  output dma_dout_10_;
  wire dma_dout_10_;
  output dma_dout_11_;
  wire dma_dout_11_;
  output dma_dout_12_;
  wire dma_dout_12_;
  output dma_dout_13_;
  wire dma_dout_13_;
  output dma_dout_14_;
  wire dma_dout_14_;
  output dma_dout_15_;
  wire dma_dout_15_;
  output dma_dout_1_;
  wire dma_dout_1_;
  output dma_dout_2_;
  wire dma_dout_2_;
  output dma_dout_3_;
  wire dma_dout_3_;
  output dma_dout_4_;
  wire dma_dout_4_;
  output dma_dout_5_;
  wire dma_dout_5_;
  output dma_dout_6_;
  wire dma_dout_6_;
  output dma_dout_7_;
  wire dma_dout_7_;
  output dma_dout_8_;
  wire dma_dout_8_;
  output dma_dout_9_;
  wire dma_dout_9_;
  input dma_en;
  wire dma_en;
  input dma_priority;
  wire dma_priority;
  output dma_ready;
  wire dma_ready;
  output dma_resp;
  wire dma_resp;
  input dma_we_0_;
  wire dma_we_0_;
  input dma_we_1_;
  wire dma_we_1_;
  input dma_wkup;
  wire dma_wkup;
  output dmem_addr_0_;
  wire dmem_addr_0_;
  output dmem_addr_10_;
  wire dmem_addr_10_;
  output dmem_addr_11_;
  wire dmem_addr_11_;
  output dmem_addr_12_;
  wire dmem_addr_12_;
  output dmem_addr_1_;
  wire dmem_addr_1_;
  output dmem_addr_2_;
  wire dmem_addr_2_;
  output dmem_addr_3_;
  wire dmem_addr_3_;
  output dmem_addr_4_;
  wire dmem_addr_4_;
  output dmem_addr_5_;
  wire dmem_addr_5_;
  output dmem_addr_6_;
  wire dmem_addr_6_;
  output dmem_addr_7_;
  wire dmem_addr_7_;
  output dmem_addr_8_;
  wire dmem_addr_8_;
  output dmem_addr_9_;
  wire dmem_addr_9_;
  output dmem_cen;
  wire dmem_cen;
  output dmem_din_0_;
  wire dmem_din_0_;
  output dmem_din_10_;
  wire dmem_din_10_;
  output dmem_din_11_;
  wire dmem_din_11_;
  output dmem_din_12_;
  wire dmem_din_12_;
  output dmem_din_13_;
  wire dmem_din_13_;
  output dmem_din_14_;
  wire dmem_din_14_;
  output dmem_din_15_;
  wire dmem_din_15_;
  output dmem_din_1_;
  wire dmem_din_1_;
  output dmem_din_2_;
  wire dmem_din_2_;
  output dmem_din_3_;
  wire dmem_din_3_;
  output dmem_din_4_;
  wire dmem_din_4_;
  output dmem_din_5_;
  wire dmem_din_5_;
  output dmem_din_6_;
  wire dmem_din_6_;
  output dmem_din_7_;
  wire dmem_din_7_;
  output dmem_din_8_;
  wire dmem_din_8_;
  output dmem_din_9_;
  wire dmem_din_9_;
  input dmem_dout_0_;
  wire dmem_dout_0_;
  input dmem_dout_10_;
  wire dmem_dout_10_;
  input dmem_dout_11_;
  wire dmem_dout_11_;
  input dmem_dout_12_;
  wire dmem_dout_12_;
  input dmem_dout_13_;
  wire dmem_dout_13_;
  input dmem_dout_14_;
  wire dmem_dout_14_;
  input dmem_dout_15_;
  wire dmem_dout_15_;
  input dmem_dout_1_;
  wire dmem_dout_1_;
  input dmem_dout_2_;
  wire dmem_dout_2_;
  input dmem_dout_3_;
  wire dmem_dout_3_;
  input dmem_dout_4_;
  wire dmem_dout_4_;
  input dmem_dout_5_;
  wire dmem_dout_5_;
  input dmem_dout_6_;
  wire dmem_dout_6_;
  input dmem_dout_7_;
  wire dmem_dout_7_;
  input dmem_dout_8_;
  wire dmem_dout_8_;
  input dmem_dout_9_;
  wire dmem_dout_9_;
  output dmem_wen_0_;
  wire dmem_wen_0_;
  output dmem_wen_1_;
  wire dmem_wen_1_;
  wire  execution_unit_0.UNUSED_inst_ad_idx ;
  wire  execution_unit_0.UNUSED_inst_ad_symb ;
  wire  execution_unit_0.alu_0.N ;
  wire  execution_unit_0.alu_0.UNUSED_inst_alu ;
  wire  execution_unit_0.alu_0.UNUSED_inst_so_call ;
  wire  execution_unit_0.alu_0.UNUSED_inst_so_push ;
  wire  execution_unit_0.alu_0.UNUSED_inst_so_reti ;
  wire  execution_unit_0.alu_0.Z ;
  wire  execution_unit_0.alu_0.alu_out_0_ ;
  wire  execution_unit_0.alu_0.alu_out_10_ ;
  wire  execution_unit_0.alu_0.alu_out_11_ ;
  wire  execution_unit_0.alu_0.alu_out_12_ ;
  wire  execution_unit_0.alu_0.alu_out_13_ ;
  wire  execution_unit_0.alu_0.alu_out_14_ ;
  wire  execution_unit_0.alu_0.alu_out_15_ ;
  wire  execution_unit_0.alu_0.alu_out_1_ ;
  wire  execution_unit_0.alu_0.alu_out_2_ ;
  wire  execution_unit_0.alu_0.alu_out_3_ ;
  wire  execution_unit_0.alu_0.alu_out_4_ ;
  wire  execution_unit_0.alu_0.alu_out_5_ ;
  wire  execution_unit_0.alu_0.alu_out_6_ ;
  wire  execution_unit_0.alu_0.alu_out_7_ ;
  wire  execution_unit_0.alu_0.alu_out_8_ ;
  wire  execution_unit_0.alu_0.alu_out_9_ ;
  wire  execution_unit_0.alu_0.alu_shift_0_ ;
  wire  execution_unit_0.alu_0.alu_shift_10_ ;
  wire  execution_unit_0.alu_0.alu_shift_11_ ;
  wire  execution_unit_0.alu_0.alu_shift_12_ ;
  wire  execution_unit_0.alu_0.alu_shift_13_ ;
  wire  execution_unit_0.alu_0.alu_shift_14_ ;
  wire  execution_unit_0.alu_0.alu_shift_1_ ;
  wire  execution_unit_0.alu_0.alu_shift_2_ ;
  wire  execution_unit_0.alu_0.alu_shift_3_ ;
  wire  execution_unit_0.alu_0.alu_shift_4_ ;
  wire  execution_unit_0.alu_0.alu_shift_5_ ;
  wire  execution_unit_0.alu_0.alu_shift_6_ ;
  wire  execution_unit_0.alu_0.alu_shift_8_ ;
  wire  execution_unit_0.alu_0.alu_shift_9_ ;
  wire  execution_unit_0.alu_0.alu_stat_0_ ;
  wire  execution_unit_0.alu_0.alu_stat_3_ ;
  wire  execution_unit_0.alu_0.alu_stat_wr_0_ ;
  wire  execution_unit_0.alu_0.alu_swpb_0_ ;
  wire  execution_unit_0.alu_0.alu_swpb_8_ ;
  wire  execution_unit_0.alu_0.exec_cycle ;
  wire  execution_unit_0.alu_0.inst_alu_0_ ;
  wire  execution_unit_0.alu_0.inst_alu_10_ ;
  wire  execution_unit_0.alu_0.inst_alu_1_ ;
  wire  execution_unit_0.alu_0.inst_alu_2_ ;
  wire  execution_unit_0.alu_0.inst_alu_3_ ;
  wire  execution_unit_0.alu_0.inst_alu_4_ ;
  wire  execution_unit_0.alu_0.inst_alu_5_ ;
  wire  execution_unit_0.alu_0.inst_alu_6_ ;
  wire  execution_unit_0.alu_0.inst_alu_7_ ;
  wire  execution_unit_0.alu_0.inst_alu_8_ ;
  wire  execution_unit_0.alu_0.inst_alu_9_ ;
  wire  execution_unit_0.alu_0.inst_bw ;
  wire  execution_unit_0.alu_0.inst_jmp_0_ ;
  wire  execution_unit_0.alu_0.inst_jmp_1_ ;
  wire  execution_unit_0.alu_0.inst_jmp_2_ ;
  wire  execution_unit_0.alu_0.inst_jmp_3_ ;
  wire  execution_unit_0.alu_0.inst_jmp_4_ ;
  wire  execution_unit_0.alu_0.inst_jmp_5_ ;
  wire  execution_unit_0.alu_0.inst_jmp_6_ ;
  wire  execution_unit_0.alu_0.inst_so_0_ ;
  wire  execution_unit_0.alu_0.inst_so_1_ ;
  wire  execution_unit_0.alu_0.inst_so_3_ ;
  wire  execution_unit_0.alu_0.inst_so_7_ ;
  wire  execution_unit_0.alu_0.op_dst_0_ ;
  wire  execution_unit_0.alu_0.op_dst_10_ ;
  wire  execution_unit_0.alu_0.op_dst_11_ ;
  wire  execution_unit_0.alu_0.op_dst_12_ ;
  wire  execution_unit_0.alu_0.op_dst_13_ ;
  wire  execution_unit_0.alu_0.op_dst_14_ ;
  wire  execution_unit_0.alu_0.op_dst_15_ ;
  wire  execution_unit_0.alu_0.op_dst_1_ ;
  wire  execution_unit_0.alu_0.op_dst_2_ ;
  wire  execution_unit_0.alu_0.op_dst_3_ ;
  wire  execution_unit_0.alu_0.op_dst_4_ ;
  wire  execution_unit_0.alu_0.op_dst_5_ ;
  wire  execution_unit_0.alu_0.op_dst_6_ ;
  wire  execution_unit_0.alu_0.op_dst_7_ ;
  wire  execution_unit_0.alu_0.op_dst_8_ ;
  wire  execution_unit_0.alu_0.op_dst_9_ ;
  wire  execution_unit_0.alu_0.status_0_ ;
  wire  execution_unit_0.alu_0.status_1_ ;
  wire  execution_unit_0.alu_0.status_2_ ;
  wire  execution_unit_0.alu_0.status_3_ ;
  wire  execution_unit_0.e_state_0_ ;
  wire  execution_unit_0.e_state_1_ ;
  wire  execution_unit_0.e_state_2_ ;
  wire  execution_unit_0.e_state_3_ ;
  wire  execution_unit_0.exec_done ;
  wire  execution_unit_0.gie ;
  wire  execution_unit_0.inst_ad_0_ ;
  wire  execution_unit_0.inst_ad_6_ ;
  wire  execution_unit_0.inst_as_0_ ;
  wire  execution_unit_0.inst_as_1_ ;
  wire  execution_unit_0.inst_as_2_ ;
  wire  execution_unit_0.inst_as_3_ ;
  wire  execution_unit_0.inst_as_4_ ;
  wire  execution_unit_0.inst_as_5_ ;
  wire  execution_unit_0.inst_as_6_ ;
  wire  execution_unit_0.inst_as_7_ ;
  wire  execution_unit_0.inst_dest_0_ ;
  wire  execution_unit_0.inst_dest_10_ ;
  wire  execution_unit_0.inst_dest_11_ ;
  wire  execution_unit_0.inst_dest_12_ ;
  wire  execution_unit_0.inst_dest_13_ ;
  wire  execution_unit_0.inst_dest_14_ ;
  wire  execution_unit_0.inst_dest_15_ ;
  wire  execution_unit_0.inst_dest_1_ ;
  wire  execution_unit_0.inst_dest_2_ ;
  wire  execution_unit_0.inst_dest_3_ ;
  wire  execution_unit_0.inst_dest_4_ ;
  wire  execution_unit_0.inst_dest_5_ ;
  wire  execution_unit_0.inst_dest_6_ ;
  wire  execution_unit_0.inst_dest_7_ ;
  wire  execution_unit_0.inst_dest_8_ ;
  wire  execution_unit_0.inst_dest_9_ ;
  wire  execution_unit_0.inst_dext_0_ ;
  wire  execution_unit_0.inst_dext_10_ ;
  wire  execution_unit_0.inst_dext_11_ ;
  wire  execution_unit_0.inst_dext_12_ ;
  wire  execution_unit_0.inst_dext_13_ ;
  wire  execution_unit_0.inst_dext_14_ ;
  wire  execution_unit_0.inst_dext_15_ ;
  wire  execution_unit_0.inst_dext_1_ ;
  wire  execution_unit_0.inst_dext_2_ ;
  wire  execution_unit_0.inst_dext_3_ ;
  wire  execution_unit_0.inst_dext_4_ ;
  wire  execution_unit_0.inst_dext_5_ ;
  wire  execution_unit_0.inst_dext_6_ ;
  wire  execution_unit_0.inst_dext_7_ ;
  wire  execution_unit_0.inst_dext_8_ ;
  wire  execution_unit_0.inst_dext_9_ ;
  wire  execution_unit_0.inst_irq_rst ;
  wire  execution_unit_0.inst_mov ;
  wire  execution_unit_0.inst_sext_0_ ;
  wire  execution_unit_0.inst_sext_10_ ;
  wire  execution_unit_0.inst_sext_11_ ;
  wire  execution_unit_0.inst_sext_12_ ;
  wire  execution_unit_0.inst_sext_13_ ;
  wire  execution_unit_0.inst_sext_14_ ;
  wire  execution_unit_0.inst_sext_15_ ;
  wire  execution_unit_0.inst_sext_1_ ;
  wire  execution_unit_0.inst_sext_2_ ;
  wire  execution_unit_0.inst_sext_3_ ;
  wire  execution_unit_0.inst_sext_4_ ;
  wire  execution_unit_0.inst_sext_5_ ;
  wire  execution_unit_0.inst_sext_6_ ;
  wire  execution_unit_0.inst_sext_7_ ;
  wire  execution_unit_0.inst_sext_8_ ;
  wire  execution_unit_0.inst_sext_9_ ;
  wire  execution_unit_0.inst_src_0_ ;
  wire  execution_unit_0.inst_src_10_ ;
  wire  execution_unit_0.inst_src_11_ ;
  wire  execution_unit_0.inst_src_12_ ;
  wire  execution_unit_0.inst_src_13_ ;
  wire  execution_unit_0.inst_src_14_ ;
  wire  execution_unit_0.inst_src_15_ ;
  wire  execution_unit_0.inst_src_1_ ;
  wire  execution_unit_0.inst_src_2_ ;
  wire  execution_unit_0.inst_src_3_ ;
  wire  execution_unit_0.inst_src_4_ ;
  wire  execution_unit_0.inst_src_5_ ;
  wire  execution_unit_0.inst_src_6_ ;
  wire  execution_unit_0.inst_src_7_ ;
  wire  execution_unit_0.inst_src_8_ ;
  wire  execution_unit_0.inst_src_9_ ;
  wire  execution_unit_0.inst_type_0_ ;
  wire  execution_unit_0.inst_type_1_ ;
  wire  execution_unit_0.inst_type_2_ ;
  wire  execution_unit_0.mab_lsb ;
  wire  execution_unit_0.mdb_in_0_ ;
  wire  execution_unit_0.mdb_in_10_ ;
  wire  execution_unit_0.mdb_in_11_ ;
  wire  execution_unit_0.mdb_in_12_ ;
  wire  execution_unit_0.mdb_in_13_ ;
  wire  execution_unit_0.mdb_in_14_ ;
  wire  execution_unit_0.mdb_in_15_ ;
  wire  execution_unit_0.mdb_in_1_ ;
  wire  execution_unit_0.mdb_in_2_ ;
  wire  execution_unit_0.mdb_in_3_ ;
  wire  execution_unit_0.mdb_in_4_ ;
  wire  execution_unit_0.mdb_in_5_ ;
  wire  execution_unit_0.mdb_in_6_ ;
  wire  execution_unit_0.mdb_in_7_ ;
  wire  execution_unit_0.mdb_in_8_ ;
  wire  execution_unit_0.mdb_in_9_ ;
  wire  execution_unit_0.mdb_in_buf_0_ ;
  wire  execution_unit_0.mdb_in_buf_10_ ;
  wire  execution_unit_0.mdb_in_buf_11_ ;
  wire  execution_unit_0.mdb_in_buf_12_ ;
  wire  execution_unit_0.mdb_in_buf_13_ ;
  wire  execution_unit_0.mdb_in_buf_14_ ;
  wire  execution_unit_0.mdb_in_buf_15_ ;
  wire  execution_unit_0.mdb_in_buf_1_ ;
  wire  execution_unit_0.mdb_in_buf_2_ ;
  wire  execution_unit_0.mdb_in_buf_3_ ;
  wire  execution_unit_0.mdb_in_buf_4_ ;
  wire  execution_unit_0.mdb_in_buf_5_ ;
  wire  execution_unit_0.mdb_in_buf_6_ ;
  wire  execution_unit_0.mdb_in_buf_7_ ;
  wire  execution_unit_0.mdb_in_buf_8_ ;
  wire  execution_unit_0.mdb_in_buf_9_ ;
  wire  execution_unit_0.mdb_in_buf_en ;
  wire  execution_unit_0.mdb_in_buf_valid ;
  wire  execution_unit_0.mdb_out_0_ ;
  wire  execution_unit_0.mdb_out_10_ ;
  wire  execution_unit_0.mdb_out_11_ ;
  wire  execution_unit_0.mdb_out_12_ ;
  wire  execution_unit_0.mdb_out_13_ ;
  wire  execution_unit_0.mdb_out_14_ ;
  wire  execution_unit_0.mdb_out_15_ ;
  wire  execution_unit_0.mdb_out_1_ ;
  wire  execution_unit_0.mdb_out_2_ ;
  wire  execution_unit_0.mdb_out_3_ ;
  wire  execution_unit_0.mdb_out_4_ ;
  wire  execution_unit_0.mdb_out_5_ ;
  wire  execution_unit_0.mdb_out_6_ ;
  wire  execution_unit_0.mdb_out_7_ ;
  wire  execution_unit_0.mdb_out_8_ ;
  wire  execution_unit_0.mdb_out_9_ ;
  wire  execution_unit_0.mdb_out_nxt_10_ ;
  wire  execution_unit_0.mdb_out_nxt_11_ ;
  wire  execution_unit_0.mdb_out_nxt_12_ ;
  wire  execution_unit_0.mdb_out_nxt_13_ ;
  wire  execution_unit_0.mdb_out_nxt_14_ ;
  wire  execution_unit_0.mdb_out_nxt_15_ ;
  wire  execution_unit_0.mdb_out_nxt_8_ ;
  wire  execution_unit_0.mdb_out_nxt_9_ ;
  wire  execution_unit_0.pc_nxt_0_ ;
  wire  execution_unit_0.pc_nxt_10_ ;
  wire  execution_unit_0.pc_nxt_11_ ;
  wire  execution_unit_0.pc_nxt_12_ ;
  wire  execution_unit_0.pc_nxt_13_ ;
  wire  execution_unit_0.pc_nxt_14_ ;
  wire  execution_unit_0.pc_nxt_15_ ;
  wire  execution_unit_0.pc_nxt_1_ ;
  wire  execution_unit_0.pc_nxt_2_ ;
  wire  execution_unit_0.pc_nxt_3_ ;
  wire  execution_unit_0.pc_nxt_4_ ;
  wire  execution_unit_0.pc_nxt_5_ ;
  wire  execution_unit_0.pc_nxt_6_ ;
  wire  execution_unit_0.pc_nxt_7_ ;
  wire  execution_unit_0.pc_nxt_8_ ;
  wire  execution_unit_0.pc_nxt_9_ ;
  wire  execution_unit_0.pc_sw_10_ ;
  wire  execution_unit_0.pc_sw_11_ ;
  wire  execution_unit_0.pc_sw_12_ ;
  wire  execution_unit_0.pc_sw_13_ ;
  wire  execution_unit_0.pc_sw_14_ ;
  wire  execution_unit_0.pc_sw_15_ ;
  wire  execution_unit_0.pc_sw_8_ ;
  wire  execution_unit_0.pc_sw_9_ ;
  wire  execution_unit_0.pc_sw_wr ;
  wire  execution_unit_0.reg_dest_wr ;
  wire  execution_unit_0.reg_incr ;
  wire  execution_unit_0.reg_pc_call ;
  wire  execution_unit_0.reg_sp_wr ;
  wire  execution_unit_0.reg_sr_clr ;
  wire  execution_unit_0.reg_sr_wr ;
  wire  execution_unit_0.reg_src_0_ ;
  wire  execution_unit_0.reg_src_10_ ;
  wire  execution_unit_0.reg_src_11_ ;
  wire  execution_unit_0.reg_src_12_ ;
  wire  execution_unit_0.reg_src_13_ ;
  wire  execution_unit_0.reg_src_14_ ;
  wire  execution_unit_0.reg_src_15_ ;
  wire  execution_unit_0.reg_src_1_ ;
  wire  execution_unit_0.reg_src_2_ ;
  wire  execution_unit_0.reg_src_3_ ;
  wire  execution_unit_0.reg_src_4_ ;
  wire  execution_unit_0.reg_src_5_ ;
  wire  execution_unit_0.reg_src_6_ ;
  wire  execution_unit_0.reg_src_7_ ;
  wire  execution_unit_0.reg_src_8_ ;
  wire  execution_unit_0.reg_src_9_ ;
  wire  execution_unit_0.register_file_0.r10_0_ ;
  wire  execution_unit_0.register_file_0.r10_10_ ;
  wire  execution_unit_0.register_file_0.r10_11_ ;
  wire  execution_unit_0.register_file_0.r10_12_ ;
  wire  execution_unit_0.register_file_0.r10_13_ ;
  wire  execution_unit_0.register_file_0.r10_14_ ;
  wire  execution_unit_0.register_file_0.r10_15_ ;
  wire  execution_unit_0.register_file_0.r10_1_ ;
  wire  execution_unit_0.register_file_0.r10_2_ ;
  wire  execution_unit_0.register_file_0.r10_3_ ;
  wire  execution_unit_0.register_file_0.r10_4_ ;
  wire  execution_unit_0.register_file_0.r10_5_ ;
  wire  execution_unit_0.register_file_0.r10_6_ ;
  wire  execution_unit_0.register_file_0.r10_7_ ;
  wire  execution_unit_0.register_file_0.r10_8_ ;
  wire  execution_unit_0.register_file_0.r10_9_ ;
  wire  execution_unit_0.register_file_0.r11_0_ ;
  wire  execution_unit_0.register_file_0.r11_10_ ;
  wire  execution_unit_0.register_file_0.r11_11_ ;
  wire  execution_unit_0.register_file_0.r11_12_ ;
  wire  execution_unit_0.register_file_0.r11_13_ ;
  wire  execution_unit_0.register_file_0.r11_14_ ;
  wire  execution_unit_0.register_file_0.r11_15_ ;
  wire  execution_unit_0.register_file_0.r11_1_ ;
  wire  execution_unit_0.register_file_0.r11_2_ ;
  wire  execution_unit_0.register_file_0.r11_3_ ;
  wire  execution_unit_0.register_file_0.r11_4_ ;
  wire  execution_unit_0.register_file_0.r11_5_ ;
  wire  execution_unit_0.register_file_0.r11_6_ ;
  wire  execution_unit_0.register_file_0.r11_7_ ;
  wire  execution_unit_0.register_file_0.r11_8_ ;
  wire  execution_unit_0.register_file_0.r11_9_ ;
  wire  execution_unit_0.register_file_0.r12_0_ ;
  wire  execution_unit_0.register_file_0.r12_10_ ;
  wire  execution_unit_0.register_file_0.r12_11_ ;
  wire  execution_unit_0.register_file_0.r12_12_ ;
  wire  execution_unit_0.register_file_0.r12_13_ ;
  wire  execution_unit_0.register_file_0.r12_14_ ;
  wire  execution_unit_0.register_file_0.r12_15_ ;
  wire  execution_unit_0.register_file_0.r12_1_ ;
  wire  execution_unit_0.register_file_0.r12_2_ ;
  wire  execution_unit_0.register_file_0.r12_3_ ;
  wire  execution_unit_0.register_file_0.r12_4_ ;
  wire  execution_unit_0.register_file_0.r12_5_ ;
  wire  execution_unit_0.register_file_0.r12_6_ ;
  wire  execution_unit_0.register_file_0.r12_7_ ;
  wire  execution_unit_0.register_file_0.r12_8_ ;
  wire  execution_unit_0.register_file_0.r12_9_ ;
  wire  execution_unit_0.register_file_0.r13_0_ ;
  wire  execution_unit_0.register_file_0.r13_10_ ;
  wire  execution_unit_0.register_file_0.r13_11_ ;
  wire  execution_unit_0.register_file_0.r13_12_ ;
  wire  execution_unit_0.register_file_0.r13_13_ ;
  wire  execution_unit_0.register_file_0.r13_14_ ;
  wire  execution_unit_0.register_file_0.r13_15_ ;
  wire  execution_unit_0.register_file_0.r13_1_ ;
  wire  execution_unit_0.register_file_0.r13_2_ ;
  wire  execution_unit_0.register_file_0.r13_3_ ;
  wire  execution_unit_0.register_file_0.r13_4_ ;
  wire  execution_unit_0.register_file_0.r13_5_ ;
  wire  execution_unit_0.register_file_0.r13_6_ ;
  wire  execution_unit_0.register_file_0.r13_7_ ;
  wire  execution_unit_0.register_file_0.r13_8_ ;
  wire  execution_unit_0.register_file_0.r13_9_ ;
  wire  execution_unit_0.register_file_0.r14_0_ ;
  wire  execution_unit_0.register_file_0.r14_10_ ;
  wire  execution_unit_0.register_file_0.r14_11_ ;
  wire  execution_unit_0.register_file_0.r14_12_ ;
  wire  execution_unit_0.register_file_0.r14_13_ ;
  wire  execution_unit_0.register_file_0.r14_14_ ;
  wire  execution_unit_0.register_file_0.r14_15_ ;
  wire  execution_unit_0.register_file_0.r14_1_ ;
  wire  execution_unit_0.register_file_0.r14_2_ ;
  wire  execution_unit_0.register_file_0.r14_3_ ;
  wire  execution_unit_0.register_file_0.r14_4_ ;
  wire  execution_unit_0.register_file_0.r14_5_ ;
  wire  execution_unit_0.register_file_0.r14_6_ ;
  wire  execution_unit_0.register_file_0.r14_7_ ;
  wire  execution_unit_0.register_file_0.r14_8_ ;
  wire  execution_unit_0.register_file_0.r14_9_ ;
  wire  execution_unit_0.register_file_0.r15_0_ ;
  wire  execution_unit_0.register_file_0.r15_10_ ;
  wire  execution_unit_0.register_file_0.r15_11_ ;
  wire  execution_unit_0.register_file_0.r15_12_ ;
  wire  execution_unit_0.register_file_0.r15_13_ ;
  wire  execution_unit_0.register_file_0.r15_14_ ;
  wire  execution_unit_0.register_file_0.r15_15_ ;
  wire  execution_unit_0.register_file_0.r15_1_ ;
  wire  execution_unit_0.register_file_0.r15_2_ ;
  wire  execution_unit_0.register_file_0.r15_3_ ;
  wire  execution_unit_0.register_file_0.r15_4_ ;
  wire  execution_unit_0.register_file_0.r15_5_ ;
  wire  execution_unit_0.register_file_0.r15_6_ ;
  wire  execution_unit_0.register_file_0.r15_7_ ;
  wire  execution_unit_0.register_file_0.r15_8_ ;
  wire  execution_unit_0.register_file_0.r15_9_ ;
  wire  execution_unit_0.register_file_0.r1_10_ ;
  wire  execution_unit_0.register_file_0.r1_11_ ;
  wire  execution_unit_0.register_file_0.r1_12_ ;
  wire  execution_unit_0.register_file_0.r1_13_ ;
  wire  execution_unit_0.register_file_0.r1_14_ ;
  wire  execution_unit_0.register_file_0.r1_15_ ;
  wire  execution_unit_0.register_file_0.r1_1_ ;
  wire  execution_unit_0.register_file_0.r1_2_ ;
  wire  execution_unit_0.register_file_0.r1_3_ ;
  wire  execution_unit_0.register_file_0.r1_4_ ;
  wire  execution_unit_0.register_file_0.r1_5_ ;
  wire  execution_unit_0.register_file_0.r1_6_ ;
  wire  execution_unit_0.register_file_0.r1_7_ ;
  wire  execution_unit_0.register_file_0.r1_8_ ;
  wire  execution_unit_0.register_file_0.r1_9_ ;
  wire  execution_unit_0.register_file_0.r2_4_ ;
  wire  execution_unit_0.register_file_0.r3_0_ ;
  wire  execution_unit_0.register_file_0.r3_10_ ;
  wire  execution_unit_0.register_file_0.r3_11_ ;
  wire  execution_unit_0.register_file_0.r3_12_ ;
  wire  execution_unit_0.register_file_0.r3_13_ ;
  wire  execution_unit_0.register_file_0.r3_14_ ;
  wire  execution_unit_0.register_file_0.r3_15_ ;
  wire  execution_unit_0.register_file_0.r3_1_ ;
  wire  execution_unit_0.register_file_0.r3_2_ ;
  wire  execution_unit_0.register_file_0.r3_3_ ;
  wire  execution_unit_0.register_file_0.r3_4_ ;
  wire  execution_unit_0.register_file_0.r3_5_ ;
  wire  execution_unit_0.register_file_0.r3_6_ ;
  wire  execution_unit_0.register_file_0.r3_7_ ;
  wire  execution_unit_0.register_file_0.r3_8_ ;
  wire  execution_unit_0.register_file_0.r3_9_ ;
  wire  execution_unit_0.register_file_0.r4_0_ ;
  wire  execution_unit_0.register_file_0.r4_10_ ;
  wire  execution_unit_0.register_file_0.r4_11_ ;
  wire  execution_unit_0.register_file_0.r4_12_ ;
  wire  execution_unit_0.register_file_0.r4_13_ ;
  wire  execution_unit_0.register_file_0.r4_14_ ;
  wire  execution_unit_0.register_file_0.r4_15_ ;
  wire  execution_unit_0.register_file_0.r4_1_ ;
  wire  execution_unit_0.register_file_0.r4_2_ ;
  wire  execution_unit_0.register_file_0.r4_3_ ;
  wire  execution_unit_0.register_file_0.r4_4_ ;
  wire  execution_unit_0.register_file_0.r4_5_ ;
  wire  execution_unit_0.register_file_0.r4_6_ ;
  wire  execution_unit_0.register_file_0.r4_7_ ;
  wire  execution_unit_0.register_file_0.r4_8_ ;
  wire  execution_unit_0.register_file_0.r4_9_ ;
  wire  execution_unit_0.register_file_0.r5_0_ ;
  wire  execution_unit_0.register_file_0.r5_10_ ;
  wire  execution_unit_0.register_file_0.r5_11_ ;
  wire  execution_unit_0.register_file_0.r5_12_ ;
  wire  execution_unit_0.register_file_0.r5_13_ ;
  wire  execution_unit_0.register_file_0.r5_14_ ;
  wire  execution_unit_0.register_file_0.r5_15_ ;
  wire  execution_unit_0.register_file_0.r5_1_ ;
  wire  execution_unit_0.register_file_0.r5_2_ ;
  wire  execution_unit_0.register_file_0.r5_3_ ;
  wire  execution_unit_0.register_file_0.r5_4_ ;
  wire  execution_unit_0.register_file_0.r5_5_ ;
  wire  execution_unit_0.register_file_0.r5_6_ ;
  wire  execution_unit_0.register_file_0.r5_7_ ;
  wire  execution_unit_0.register_file_0.r5_8_ ;
  wire  execution_unit_0.register_file_0.r5_9_ ;
  wire  execution_unit_0.register_file_0.r6_0_ ;
  wire  execution_unit_0.register_file_0.r6_10_ ;
  wire  execution_unit_0.register_file_0.r6_11_ ;
  wire  execution_unit_0.register_file_0.r6_12_ ;
  wire  execution_unit_0.register_file_0.r6_13_ ;
  wire  execution_unit_0.register_file_0.r6_14_ ;
  wire  execution_unit_0.register_file_0.r6_15_ ;
  wire  execution_unit_0.register_file_0.r6_1_ ;
  wire  execution_unit_0.register_file_0.r6_2_ ;
  wire  execution_unit_0.register_file_0.r6_3_ ;
  wire  execution_unit_0.register_file_0.r6_4_ ;
  wire  execution_unit_0.register_file_0.r6_5_ ;
  wire  execution_unit_0.register_file_0.r6_6_ ;
  wire  execution_unit_0.register_file_0.r6_7_ ;
  wire  execution_unit_0.register_file_0.r6_8_ ;
  wire  execution_unit_0.register_file_0.r6_9_ ;
  wire  execution_unit_0.register_file_0.r7_0_ ;
  wire  execution_unit_0.register_file_0.r7_10_ ;
  wire  execution_unit_0.register_file_0.r7_11_ ;
  wire  execution_unit_0.register_file_0.r7_12_ ;
  wire  execution_unit_0.register_file_0.r7_13_ ;
  wire  execution_unit_0.register_file_0.r7_14_ ;
  wire  execution_unit_0.register_file_0.r7_15_ ;
  wire  execution_unit_0.register_file_0.r7_1_ ;
  wire  execution_unit_0.register_file_0.r7_2_ ;
  wire  execution_unit_0.register_file_0.r7_3_ ;
  wire  execution_unit_0.register_file_0.r7_4_ ;
  wire  execution_unit_0.register_file_0.r7_5_ ;
  wire  execution_unit_0.register_file_0.r7_6_ ;
  wire  execution_unit_0.register_file_0.r7_7_ ;
  wire  execution_unit_0.register_file_0.r7_8_ ;
  wire  execution_unit_0.register_file_0.r7_9_ ;
  wire  execution_unit_0.register_file_0.r8_0_ ;
  wire  execution_unit_0.register_file_0.r8_10_ ;
  wire  execution_unit_0.register_file_0.r8_11_ ;
  wire  execution_unit_0.register_file_0.r8_12_ ;
  wire  execution_unit_0.register_file_0.r8_13_ ;
  wire  execution_unit_0.register_file_0.r8_14_ ;
  wire  execution_unit_0.register_file_0.r8_15_ ;
  wire  execution_unit_0.register_file_0.r8_1_ ;
  wire  execution_unit_0.register_file_0.r8_2_ ;
  wire  execution_unit_0.register_file_0.r8_3_ ;
  wire  execution_unit_0.register_file_0.r8_4_ ;
  wire  execution_unit_0.register_file_0.r8_5_ ;
  wire  execution_unit_0.register_file_0.r8_6_ ;
  wire  execution_unit_0.register_file_0.r8_7_ ;
  wire  execution_unit_0.register_file_0.r8_8_ ;
  wire  execution_unit_0.register_file_0.r8_9_ ;
  wire  execution_unit_0.register_file_0.r9_0_ ;
  wire  execution_unit_0.register_file_0.r9_10_ ;
  wire  execution_unit_0.register_file_0.r9_11_ ;
  wire  execution_unit_0.register_file_0.r9_12_ ;
  wire  execution_unit_0.register_file_0.r9_13_ ;
  wire  execution_unit_0.register_file_0.r9_14_ ;
  wire  execution_unit_0.register_file_0.r9_15_ ;
  wire  execution_unit_0.register_file_0.r9_1_ ;
  wire  execution_unit_0.register_file_0.r9_2_ ;
  wire  execution_unit_0.register_file_0.r9_3_ ;
  wire  execution_unit_0.register_file_0.r9_4_ ;
  wire  execution_unit_0.register_file_0.r9_5_ ;
  wire  execution_unit_0.register_file_0.r9_6_ ;
  wire  execution_unit_0.register_file_0.r9_7_ ;
  wire  execution_unit_0.register_file_0.r9_8_ ;
  wire  execution_unit_0.register_file_0.r9_9_ ;
  wire  frontend_0.e_state_nxt_0_ ;
  wire  frontend_0.e_state_nxt_1_ ;
  wire  frontend_0.e_state_nxt_2_ ;
  wire  frontend_0.e_state_nxt_3_ ;
  wire  frontend_0.exec_dext_rdy ;
  wire  frontend_0.exec_dst_wr ;
  wire  frontend_0.exec_jmp ;
  wire  frontend_0.exec_src_wr ;
  wire  frontend_0.fe_pmem_wait ;
  wire  frontend_0.i_state_0_ ;
  wire  frontend_0.i_state_1_ ;
  wire  frontend_0.i_state_2_ ;
  wire  frontend_0.i_state_nxt_0_ ;
  wire  frontend_0.i_state_nxt_1_ ;
  wire  frontend_0.i_state_nxt_2_ ;
  wire  frontend_0.inst_dest_bin_0_ ;
  wire  frontend_0.inst_dest_bin_1_ ;
  wire  frontend_0.inst_dest_bin_2_ ;
  wire  frontend_0.inst_dest_bin_3_ ;
  wire  frontend_0.inst_jmp_bin_0_ ;
  wire  frontend_0.inst_jmp_bin_1_ ;
  wire  frontend_0.inst_jmp_bin_2_ ;
  wire  frontend_0.inst_src_bin_0_ ;
  wire  frontend_0.inst_src_bin_1_ ;
  wire  frontend_0.inst_sz_0_ ;
  wire  frontend_0.inst_sz_1_ ;
  wire  frontend_0.irq_addr_1_ ;
  wire  frontend_0.irq_addr_2_ ;
  wire  frontend_0.irq_addr_3_ ;
  wire  frontend_0.irq_addr_4_ ;
  wire  frontend_0.mb_en ;
  wire  frontend_0.pmem_busy ;
  wire  frontend_0.wdt_irq ;
  input irq_0_;
  wire irq_0_;
  input irq_10_;
  wire irq_10_;
  input irq_11_;
  wire irq_11_;
  input irq_12_;
  wire irq_12_;
  input irq_13_;
  wire irq_13_;
  input irq_1_;
  wire irq_1_;
  input irq_2_;
  wire irq_2_;
  input irq_3_;
  wire irq_3_;
  input irq_4_;
  wire irq_4_;
  input irq_5_;
  wire irq_5_;
  input irq_6_;
  wire irq_6_;
  input irq_7_;
  wire irq_7_;
  input irq_8_;
  wire irq_8_;
  input irq_9_;
  wire irq_9_;
  output irq_acc_0_;
  wire irq_acc_0_;
  output irq_acc_10_;
  wire irq_acc_10_;
  output irq_acc_11_;
  wire irq_acc_11_;
  output irq_acc_12_;
  wire irq_acc_12_;
  output irq_acc_13_;
  wire irq_acc_13_;
  output irq_acc_1_;
  wire irq_acc_1_;
  output irq_acc_2_;
  wire irq_acc_2_;
  output irq_acc_3_;
  wire irq_acc_3_;
  output irq_acc_4_;
  wire irq_acc_4_;
  output irq_acc_5_;
  wire irq_acc_5_;
  output irq_acc_6_;
  wire irq_acc_6_;
  output irq_acc_7_;
  wire irq_acc_7_;
  output irq_acc_8_;
  wire irq_acc_8_;
  output irq_acc_9_;
  wire irq_acc_9_;
  input lfxt_clk;
  wire lfxt_clk;
  output lfxt_enable;
  wire lfxt_enable;
  output lfxt_wkup;
  wire lfxt_wkup;
  output mclk;
  wire mclk;
  wire  mem_backbone_0.eu_mdb_in_sel_0_ ;
  wire  mem_backbone_0.eu_mdb_in_sel_1_ ;
  wire  mem_backbone_0.eu_per_en ;
  wire  mem_backbone_0.eu_pmem_en ;
  wire  mem_backbone_0.ext_mem_din_sel ;
  wire  mem_backbone_0.ext_per_en ;
  wire  mem_backbone_0.ext_pmem_en ;
  wire  mem_backbone_0.fe_pmem_en ;
  wire  mem_backbone_0.fe_pmem_en_dly ;
  wire  mem_backbone_0.per_dout_0_ ;
  wire  mem_backbone_0.per_dout_10_ ;
  wire  mem_backbone_0.per_dout_11_ ;
  wire  mem_backbone_0.per_dout_12_ ;
  wire  mem_backbone_0.per_dout_13_ ;
  wire  mem_backbone_0.per_dout_14_ ;
  wire  mem_backbone_0.per_dout_15_ ;
  wire  mem_backbone_0.per_dout_1_ ;
  wire  mem_backbone_0.per_dout_2_ ;
  wire  mem_backbone_0.per_dout_3_ ;
  wire  mem_backbone_0.per_dout_4_ ;
  wire  mem_backbone_0.per_dout_5_ ;
  wire  mem_backbone_0.per_dout_6_ ;
  wire  mem_backbone_0.per_dout_7_ ;
  wire  mem_backbone_0.per_dout_8_ ;
  wire  mem_backbone_0.per_dout_9_ ;
  wire  mem_backbone_0.per_dout_val_0_ ;
  wire  mem_backbone_0.per_dout_val_10_ ;
  wire  mem_backbone_0.per_dout_val_11_ ;
  wire  mem_backbone_0.per_dout_val_12_ ;
  wire  mem_backbone_0.per_dout_val_13_ ;
  wire  mem_backbone_0.per_dout_val_14_ ;
  wire  mem_backbone_0.per_dout_val_15_ ;
  wire  mem_backbone_0.per_dout_val_1_ ;
  wire  mem_backbone_0.per_dout_val_2_ ;
  wire  mem_backbone_0.per_dout_val_3_ ;
  wire  mem_backbone_0.per_dout_val_4_ ;
  wire  mem_backbone_0.per_dout_val_5_ ;
  wire  mem_backbone_0.per_dout_val_6_ ;
  wire  mem_backbone_0.per_dout_val_7_ ;
  wire  mem_backbone_0.per_dout_val_8_ ;
  wire  mem_backbone_0.per_dout_val_9_ ;
  wire  mem_backbone_0.pmem_dout_bckup_0_ ;
  wire  mem_backbone_0.pmem_dout_bckup_10_ ;
  wire  mem_backbone_0.pmem_dout_bckup_11_ ;
  wire  mem_backbone_0.pmem_dout_bckup_12_ ;
  wire  mem_backbone_0.pmem_dout_bckup_13_ ;
  wire  mem_backbone_0.pmem_dout_bckup_14_ ;
  wire  mem_backbone_0.pmem_dout_bckup_15_ ;
  wire  mem_backbone_0.pmem_dout_bckup_1_ ;
  wire  mem_backbone_0.pmem_dout_bckup_2_ ;
  wire  mem_backbone_0.pmem_dout_bckup_3_ ;
  wire  mem_backbone_0.pmem_dout_bckup_4_ ;
  wire  mem_backbone_0.pmem_dout_bckup_5_ ;
  wire  mem_backbone_0.pmem_dout_bckup_6_ ;
  wire  mem_backbone_0.pmem_dout_bckup_7_ ;
  wire  mem_backbone_0.pmem_dout_bckup_8_ ;
  wire  mem_backbone_0.pmem_dout_bckup_9_ ;
  wire  mem_backbone_0.pmem_dout_bckup_sel ;
  wire  multiplier_0.acc_sel ;
  wire  multiplier_0.cycle_0_ ;
  wire  multiplier_0.cycle_1_ ;
  wire  multiplier_0.op1_0_ ;
  wire  multiplier_0.op1_10_ ;
  wire  multiplier_0.op1_11_ ;
  wire  multiplier_0.op1_12_ ;
  wire  multiplier_0.op1_13_ ;
  wire  multiplier_0.op1_14_ ;
  wire  multiplier_0.op1_15_ ;
  wire  multiplier_0.op1_1_ ;
  wire  multiplier_0.op1_2_ ;
  wire  multiplier_0.op1_3_ ;
  wire  multiplier_0.op1_4_ ;
  wire  multiplier_0.op1_5_ ;
  wire  multiplier_0.op1_6_ ;
  wire  multiplier_0.op1_7_ ;
  wire  multiplier_0.op1_8_ ;
  wire  multiplier_0.op1_9_ ;
  wire  multiplier_0.op2_0_ ;
  wire  multiplier_0.op2_10_ ;
  wire  multiplier_0.op2_11_ ;
  wire  multiplier_0.op2_12_ ;
  wire  multiplier_0.op2_13_ ;
  wire  multiplier_0.op2_14_ ;
  wire  multiplier_0.op2_15_ ;
  wire  multiplier_0.op2_1_ ;
  wire  multiplier_0.op2_2_ ;
  wire  multiplier_0.op2_3_ ;
  wire  multiplier_0.op2_4_ ;
  wire  multiplier_0.op2_5_ ;
  wire  multiplier_0.op2_6_ ;
  wire  multiplier_0.op2_7_ ;
  wire  multiplier_0.op2_8_ ;
  wire  multiplier_0.op2_9_ ;
  wire  multiplier_0.op2_wr ;
  wire  multiplier_0.per_dout_0_ ;
  wire  multiplier_0.per_dout_10_ ;
  wire  multiplier_0.per_dout_11_ ;
  wire  multiplier_0.per_dout_12_ ;
  wire  multiplier_0.per_dout_13_ ;
  wire  multiplier_0.per_dout_14_ ;
  wire  multiplier_0.per_dout_15_ ;
  wire  multiplier_0.per_dout_1_ ;
  wire  multiplier_0.per_dout_2_ ;
  wire  multiplier_0.per_dout_3_ ;
  wire  multiplier_0.per_dout_4_ ;
  wire  multiplier_0.per_dout_5_ ;
  wire  multiplier_0.per_dout_6_ ;
  wire  multiplier_0.per_dout_7_ ;
  wire  multiplier_0.per_dout_8_ ;
  wire  multiplier_0.per_dout_9_ ;
  wire  multiplier_0.reshi_0_ ;
  wire  multiplier_0.reshi_10_ ;
  wire  multiplier_0.reshi_11_ ;
  wire  multiplier_0.reshi_12_ ;
  wire  multiplier_0.reshi_13_ ;
  wire  multiplier_0.reshi_14_ ;
  wire  multiplier_0.reshi_15_ ;
  wire  multiplier_0.reshi_1_ ;
  wire  multiplier_0.reshi_2_ ;
  wire  multiplier_0.reshi_3_ ;
  wire  multiplier_0.reshi_4_ ;
  wire  multiplier_0.reshi_5_ ;
  wire  multiplier_0.reshi_6_ ;
  wire  multiplier_0.reshi_7_ ;
  wire  multiplier_0.reshi_8_ ;
  wire  multiplier_0.reshi_9_ ;
  wire  multiplier_0.reslo_0_ ;
  wire  multiplier_0.reslo_10_ ;
  wire  multiplier_0.reslo_11_ ;
  wire  multiplier_0.reslo_12_ ;
  wire  multiplier_0.reslo_13_ ;
  wire  multiplier_0.reslo_14_ ;
  wire  multiplier_0.reslo_15_ ;
  wire  multiplier_0.reslo_1_ ;
  wire  multiplier_0.reslo_2_ ;
  wire  multiplier_0.reslo_3_ ;
  wire  multiplier_0.reslo_4_ ;
  wire  multiplier_0.reslo_5_ ;
  wire  multiplier_0.reslo_6_ ;
  wire  multiplier_0.reslo_7_ ;
  wire  multiplier_0.reslo_8_ ;
  wire  multiplier_0.reslo_9_ ;
  wire  multiplier_0.sign_sel ;
  wire  multiplier_0.sumext_0_ ;
  wire  multiplier_0.sumext_10_ ;
  input nmi;
  wire nmi;
  output per_addr_0_;
  wire per_addr_0_;
  output per_addr_10_;
  wire per_addr_10_;
  output per_addr_11_;
  wire per_addr_11_;
  output per_addr_12_;
  wire per_addr_12_;
  output per_addr_13_;
  wire per_addr_13_;
  output per_addr_1_;
  wire per_addr_1_;
  output per_addr_2_;
  wire per_addr_2_;
  output per_addr_3_;
  wire per_addr_3_;
  output per_addr_4_;
  wire per_addr_4_;
  output per_addr_5_;
  wire per_addr_5_;
  output per_addr_6_;
  wire per_addr_6_;
  output per_addr_7_;
  wire per_addr_7_;
  output per_addr_8_;
  wire per_addr_8_;
  output per_addr_9_;
  wire per_addr_9_;
  output per_din_0_;
  wire per_din_0_;
  output per_din_10_;
  wire per_din_10_;
  output per_din_11_;
  wire per_din_11_;
  output per_din_12_;
  wire per_din_12_;
  output per_din_13_;
  wire per_din_13_;
  output per_din_14_;
  wire per_din_14_;
  output per_din_15_;
  wire per_din_15_;
  output per_din_1_;
  wire per_din_1_;
  output per_din_2_;
  wire per_din_2_;
  output per_din_3_;
  wire per_din_3_;
  output per_din_4_;
  wire per_din_4_;
  output per_din_5_;
  wire per_din_5_;
  output per_din_6_;
  wire per_din_6_;
  output per_din_7_;
  wire per_din_7_;
  output per_din_8_;
  wire per_din_8_;
  output per_din_9_;
  wire per_din_9_;
  input per_dout_0_;
  wire per_dout_0_;
  input per_dout_10_;
  wire per_dout_10_;
  input per_dout_11_;
  wire per_dout_11_;
  input per_dout_12_;
  wire per_dout_12_;
  input per_dout_13_;
  wire per_dout_13_;
  input per_dout_14_;
  wire per_dout_14_;
  input per_dout_15_;
  wire per_dout_15_;
  input per_dout_1_;
  wire per_dout_1_;
  input per_dout_2_;
  wire per_dout_2_;
  input per_dout_3_;
  wire per_dout_3_;
  input per_dout_4_;
  wire per_dout_4_;
  input per_dout_5_;
  wire per_dout_5_;
  input per_dout_6_;
  wire per_dout_6_;
  input per_dout_7_;
  wire per_dout_7_;
  input per_dout_8_;
  wire per_dout_8_;
  input per_dout_9_;
  wire per_dout_9_;
  output per_en;
  wire per_en;
  output per_we_0_;
  wire per_we_0_;
  output per_we_1_;
  wire per_we_1_;
  output pmem_addr_0_;
  wire pmem_addr_0_;
  output pmem_addr_10_;
  wire pmem_addr_10_;
  output pmem_addr_11_;
  wire pmem_addr_11_;
  output pmem_addr_12_;
  wire pmem_addr_12_;
  output pmem_addr_13_;
  wire pmem_addr_13_;
  output pmem_addr_1_;
  wire pmem_addr_1_;
  output pmem_addr_2_;
  wire pmem_addr_2_;
  output pmem_addr_3_;
  wire pmem_addr_3_;
  output pmem_addr_4_;
  wire pmem_addr_4_;
  output pmem_addr_5_;
  wire pmem_addr_5_;
  output pmem_addr_6_;
  wire pmem_addr_6_;
  output pmem_addr_7_;
  wire pmem_addr_7_;
  output pmem_addr_8_;
  wire pmem_addr_8_;
  output pmem_addr_9_;
  wire pmem_addr_9_;
  output pmem_cen;
  wire pmem_cen;
  output pmem_din_0_;
  wire pmem_din_0_;
  output pmem_din_10_;
  wire pmem_din_10_;
  output pmem_din_11_;
  wire pmem_din_11_;
  output pmem_din_12_;
  wire pmem_din_12_;
  output pmem_din_13_;
  wire pmem_din_13_;
  output pmem_din_14_;
  wire pmem_din_14_;
  output pmem_din_15_;
  wire pmem_din_15_;
  output pmem_din_1_;
  wire pmem_din_1_;
  output pmem_din_2_;
  wire pmem_din_2_;
  output pmem_din_3_;
  wire pmem_din_3_;
  output pmem_din_4_;
  wire pmem_din_4_;
  output pmem_din_5_;
  wire pmem_din_5_;
  output pmem_din_6_;
  wire pmem_din_6_;
  output pmem_din_7_;
  wire pmem_din_7_;
  output pmem_din_8_;
  wire pmem_din_8_;
  output pmem_din_9_;
  wire pmem_din_9_;
  input pmem_dout_0_;
  wire pmem_dout_0_;
  input pmem_dout_10_;
  wire pmem_dout_10_;
  input pmem_dout_11_;
  wire pmem_dout_11_;
  input pmem_dout_12_;
  wire pmem_dout_12_;
  input pmem_dout_13_;
  wire pmem_dout_13_;
  input pmem_dout_14_;
  wire pmem_dout_14_;
  input pmem_dout_15_;
  wire pmem_dout_15_;
  input pmem_dout_1_;
  wire pmem_dout_1_;
  input pmem_dout_2_;
  wire pmem_dout_2_;
  input pmem_dout_3_;
  wire pmem_dout_3_;
  input pmem_dout_4_;
  wire pmem_dout_4_;
  input pmem_dout_5_;
  wire pmem_dout_5_;
  input pmem_dout_6_;
  wire pmem_dout_6_;
  input pmem_dout_7_;
  wire pmem_dout_7_;
  input pmem_dout_8_;
  wire pmem_dout_8_;
  input pmem_dout_9_;
  wire pmem_dout_9_;
  output pmem_wen_0_;
  wire pmem_wen_0_;
  output pmem_wen_1_;
  wire pmem_wen_1_;
  output puc_rst;
  wire puc_rst;
  input reset_n;
  wire reset_n;
  input scan_enable;
  wire scan_enable;
  input scan_mode;
  wire scan_mode;
  wire  sfr_0.cpu_nr_rd_10_ ;
  wire  sfr_0.cpu_nr_rd_11_ ;
  wire  sfr_0.cpu_nr_rd_12_ ;
  wire  sfr_0.cpu_nr_rd_13_ ;
  wire  sfr_0.cpu_nr_rd_2_ ;
  wire  sfr_0.cpu_nr_rd_3_ ;
  wire  sfr_0.cpu_nr_rd_4_ ;
  wire  sfr_0.cpu_nr_rd_5_ ;
  wire  sfr_0.cpu_nr_rd_6_ ;
  wire  sfr_0.cpu_nr_rd_7_ ;
  wire  sfr_0.cpu_nr_rd_9_ ;
  wire  sfr_0.ie1_0_ ;
  wire  sfr_0.ifg1_0_ ;
  wire  sfr_0.per_dout_0_ ;
  wire  sfr_0.per_dout_14_ ;
  wire  sfr_0.per_dout_15_ ;
  wire  sfr_0.per_dout_1_ ;
  wire  sfr_0.per_dout_8_ ;
  wire  sfr_0.wdtifg_sw_clr ;
  wire  sfr_0.wdtifg_sw_set ;
  output smclk;
  wire smclk;
  output smclk_en;
  wire smclk_en;
  wire  watchdog_0.per_dout_0_ ;
  wire  watchdog_0.per_dout_11_ ;
  wire  watchdog_0.per_dout_1_ ;
  wire  watchdog_0.per_dout_2_ ;
  wire  watchdog_0.per_dout_4_ ;
  wire  watchdog_0.per_dout_7_ ;
  wire  watchdog_0.wdtcnt_0_ ;
  wire  watchdog_0.wdtcnt_10_ ;
  wire  watchdog_0.wdtcnt_11_ ;
  wire  watchdog_0.wdtcnt_12_ ;
  wire  watchdog_0.wdtcnt_13_ ;
  wire  watchdog_0.wdtcnt_14_ ;
  wire  watchdog_0.wdtcnt_15_ ;
  wire  watchdog_0.wdtcnt_1_ ;
  wire  watchdog_0.wdtcnt_2_ ;
  wire  watchdog_0.wdtcnt_3_ ;
  wire  watchdog_0.wdtcnt_4_ ;
  wire  watchdog_0.wdtcnt_5_ ;
  wire  watchdog_0.wdtcnt_6_ ;
  wire  watchdog_0.wdtcnt_7_ ;
  wire  watchdog_0.wdtcnt_8_ ;
  wire  watchdog_0.wdtcnt_9_ ;
  wire  watchdog_0.wdtctl_0_ ;
  wire  watchdog_0.wdtctl_1_ ;
  wire  watchdog_0.wdtctl_2_ ;
  wire  watchdog_0.wdtctl_4_ ;
  wire  watchdog_0.wdtctl_7_ ;
  input wkup;
  wire wkup;
  INVX1 _05697_ (
    .A( multiplier_0.per_dout_0_ ),
    .Y(_00045_)
  );
  INVX1 _05698_ (
    .A( multiplier_0.per_dout_1_ ),
    .Y(_00046_)
  );
  INVX1 _05699_ (
    .A( multiplier_0.per_dout_2_ ),
    .Y(_00047_)
  );
  INVX1 _05700_ (
    .A( multiplier_0.per_dout_3_ ),
    .Y(_00000_)
  );
  INVX1 _05701_ (
    .A( multiplier_0.per_dout_4_ ),
    .Y(_00001_)
  );
  INVX1 _05702_ (
    .A( multiplier_0.per_dout_5_ ),
    .Y(_00002_)
  );
  INVX1 _05703_ (
    .A( multiplier_0.per_dout_6_ ),
    .Y(_00003_)
  );
  INVX1 _05704_ (
    .A( multiplier_0.per_dout_7_ ),
    .Y(_00004_)
  );
  INVX1 _05705_ (
    .A( multiplier_0.per_dout_8_ ),
    .Y(_00005_)
  );
  INVX1 _05706_ (
    .A( multiplier_0.per_dout_9_ ),
    .Y(_00006_)
  );
  INVX1 _05707_ (
    .A( multiplier_0.per_dout_10_ ),
    .Y(_00007_)
  );
  INVX1 _05708_ (
    .A( multiplier_0.per_dout_11_ ),
    .Y(_00008_)
  );
  INVX1 _05709_ (
    .A( multiplier_0.per_dout_12_ ),
    .Y(_00009_)
  );
  INVX1 _05710_ (
    .A( multiplier_0.per_dout_13_ ),
    .Y(_00010_)
  );
  INVX1 _05711_ (
    .A( multiplier_0.per_dout_14_ ),
    .Y(_00011_)
  );
  INVX1 _05712_ (
    .A( multiplier_0.per_dout_15_ ),
    .Y(_00012_)
  );
  NOR2X1 _05713_ (
    .A(1'h0),
    .B(per_dout_0_),
    .Y(_00013_)
  );
  NOR2X1 _05714_ (
    .A( sfr_0.per_dout_0_ ),
    .B( watchdog_0.per_dout_0_ ),
    .Y(_00014_)
  );
  NAND3X1 _05715_ (
    .A(_00045_),
    .B(_00013_),
    .C(_00014_),
    .Y( mem_backbone_0.per_dout_0_ )
  );
  NOR2X1 _05716_ (
    .A( clock_module_0.bcsctl2_rd_1_ ),
    .B(per_dout_1_),
    .Y(_00015_)
  );
  NOR2X1 _05717_ (
    .A( sfr_0.per_dout_1_ ),
    .B( watchdog_0.per_dout_1_ ),
    .Y(_00016_)
  );
  NAND3X1 _05718_ (
    .A(_00046_),
    .B(_00015_),
    .C(_00016_),
    .Y( mem_backbone_0.per_dout_1_ )
  );
  NOR2X1 _05719_ (
    .A( clock_module_0.bcsctl2_rd_2_ ),
    .B(per_dout_2_),
    .Y(_00017_)
  );
  NOR2X1 _05720_ (
    .A( sfr_0.cpu_nr_rd_2_ ),
    .B( watchdog_0.per_dout_2_ ),
    .Y(_00018_)
  );
  NAND3X1 _05721_ (
    .A(_00047_),
    .B(_00017_),
    .C(_00018_),
    .Y( mem_backbone_0.per_dout_2_ )
  );
  NOR2X1 _05722_ (
    .A( clock_module_0.bcsctl2_rd_3_ ),
    .B(per_dout_3_),
    .Y(_00019_)
  );
  NOR2X1 _05723_ (
    .A( sfr_0.cpu_nr_rd_3_ ),
    .B(1'h0),
    .Y(_00020_)
  );
  NAND3X1 _05724_ (
    .A(_00000_),
    .B(_00019_),
    .C(_00020_),
    .Y( mem_backbone_0.per_dout_3_ )
  );
  NOR2X1 _05725_ (
    .A(1'h0),
    .B(per_dout_4_),
    .Y(_00021_)
  );
  NOR2X1 _05726_ (
    .A( sfr_0.cpu_nr_rd_4_ ),
    .B( watchdog_0.per_dout_4_ ),
    .Y(_00022_)
  );
  NAND3X1 _05727_ (
    .A(_00001_),
    .B(_00021_),
    .C(_00022_),
    .Y( mem_backbone_0.per_dout_4_ )
  );
  NOR2X1 _05728_ (
    .A(1'h0),
    .B(per_dout_5_),
    .Y(_00023_)
  );
  NOR2X1 _05729_ (
    .A( sfr_0.cpu_nr_rd_5_ ),
    .B(1'h0),
    .Y(_00024_)
  );
  NAND3X1 _05730_ (
    .A(_00002_),
    .B(_00023_),
    .C(_00024_),
    .Y( mem_backbone_0.per_dout_5_ )
  );
  NOR2X1 _05731_ (
    .A(1'h0),
    .B(per_dout_6_),
    .Y(_00025_)
  );
  NOR2X1 _05732_ (
    .A( sfr_0.cpu_nr_rd_6_ ),
    .B(1'h0),
    .Y(_00026_)
  );
  NAND3X1 _05733_ (
    .A(_00003_),
    .B(_00025_),
    .C(_00026_),
    .Y( mem_backbone_0.per_dout_6_ )
  );
  NOR2X1 _05734_ (
    .A(1'h0),
    .B(per_dout_7_),
    .Y(_00027_)
  );
  NOR2X1 _05735_ (
    .A( sfr_0.cpu_nr_rd_7_ ),
    .B( watchdog_0.per_dout_7_ ),
    .Y(_00028_)
  );
  NAND3X1 _05736_ (
    .A(_00004_),
    .B(_00027_),
    .C(_00028_),
    .Y( mem_backbone_0.per_dout_7_ )
  );
  NOR2X1 _05737_ (
    .A(1'h0),
    .B(per_dout_8_),
    .Y(_00029_)
  );
  NOR2X1 _05738_ (
    .A( sfr_0.per_dout_8_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00030_)
  );
  NAND3X1 _05739_ (
    .A(_00005_),
    .B(_00029_),
    .C(_00030_),
    .Y( mem_backbone_0.per_dout_8_ )
  );
  NOR2X1 _05740_ (
    .A(1'h0),
    .B(per_dout_9_),
    .Y(_00031_)
  );
  NOR2X1 _05741_ (
    .A( sfr_0.cpu_nr_rd_9_ ),
    .B(1'h0),
    .Y(_00032_)
  );
  NAND3X1 _05742_ (
    .A(_00006_),
    .B(_00031_),
    .C(_00032_),
    .Y( mem_backbone_0.per_dout_9_ )
  );
  NOR2X1 _05743_ (
    .A(1'h0),
    .B(per_dout_10_),
    .Y(_00033_)
  );
  NOR2X1 _05744_ (
    .A( sfr_0.cpu_nr_rd_10_ ),
    .B(1'h0),
    .Y(_00034_)
  );
  NAND3X1 _05745_ (
    .A(_00007_),
    .B(_00033_),
    .C(_00034_),
    .Y( mem_backbone_0.per_dout_10_ )
  );
  NOR2X1 _05746_ (
    .A(1'h0),
    .B(per_dout_11_),
    .Y(_00035_)
  );
  NOR2X1 _05747_ (
    .A( sfr_0.cpu_nr_rd_11_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00036_)
  );
  NAND3X1 _05748_ (
    .A(_00008_),
    .B(_00035_),
    .C(_00036_),
    .Y( mem_backbone_0.per_dout_11_ )
  );
  NOR2X1 _05749_ (
    .A( clock_module_0.bcsctl1_rd_12_ ),
    .B(per_dout_12_),
    .Y(_00037_)
  );
  NOR2X1 _05750_ (
    .A( sfr_0.cpu_nr_rd_12_ ),
    .B(1'h0),
    .Y(_00038_)
  );
  NAND3X1 _05751_ (
    .A(_00009_),
    .B(_00037_),
    .C(_00038_),
    .Y( mem_backbone_0.per_dout_12_ )
  );
  NOR2X1 _05752_ (
    .A( clock_module_0.bcsctl1_rd_13_ ),
    .B(per_dout_13_),
    .Y(_00039_)
  );
  NOR2X1 _05753_ (
    .A( sfr_0.cpu_nr_rd_13_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00040_)
  );
  NAND3X1 _05754_ (
    .A(_00010_),
    .B(_00039_),
    .C(_00040_),
    .Y( mem_backbone_0.per_dout_13_ )
  );
  NOR2X1 _05755_ (
    .A(1'h0),
    .B(per_dout_14_),
    .Y(_00041_)
  );
  NOR2X1 _05756_ (
    .A( sfr_0.per_dout_14_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y(_00042_)
  );
  NAND3X1 _05757_ (
    .A(_00011_),
    .B(_00041_),
    .C(_00042_),
    .Y( mem_backbone_0.per_dout_14_ )
  );
  NOR2X1 _05758_ (
    .A(1'h0),
    .B(per_dout_15_),
    .Y(_00043_)
  );
  NOR2X1 _05759_ (
    .A( sfr_0.per_dout_15_ ),
    .B(1'h0),
    .Y(_00044_)
  );
  NAND3X1 _05760_ (
    .A(_00012_),
    .B(_00043_),
    .C(_00044_),
    .Y( mem_backbone_0.per_dout_15_ )
  );
  INVX1 _05761_ (
    .A( clock_module_0.aclk_div_0_ ),
    .Y(_00097_)
  );
  INVX1 _05762_ (
    .A(reset_n),
    .Y( clock_module_0.por_a )
  );
  INVX1 _05763_ (
    .A(dbg_en),
    .Y( clock_module_0.dbg_rst_nxt )
  );
  INVX1 _05764_ (
    .A( clock_module_0.puc_noscan_n ),
    .Y(_05695_)
  );
  INVX1 _05765_ (
    .A(_05637_),
    .Y(_00098_)
  );
  INVX1 _05766_ (
    .A(_05639_),
    .Y(_00099_)
  );
  INVX1 _05767_ (
    .A(_05633_),
    .Y(_00100_)
  );
  INVX1 _05768_ (
    .A( clock_module_0.bcsctl2_2_ ),
    .Y(_00101_)
  );
  INVX1 _05769_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .Y(_00102_)
  );
  INVX1 _05770_ (
    .A( clock_module_0.lfxt_clk_dly ),
    .Y(_00103_)
  );
  INVX1 _05771_ (
    .A( clock_module_0.oscoff ),
    .Y(_00104_)
  );
  INVX1 _05772_ (
    .A( clock_module_0.aclk_div_1_ ),
    .Y(_00105_)
  );
  INVX1 _05773_ (
    .A( clock_module_0.smclk_div_1_ ),
    .Y(_00106_)
  );
  INVX1 _05774_ (
    .A( clock_module_0.smclk_div_2_ ),
    .Y(_00107_)
  );
  INVX1 _05775_ (
    .A( clock_module_0.por ),
    .Y(_00050_)
  );
  NOR2X1 _05776_ (
    .A( clock_module_0.dbg_rst_nxt ),
    .B( clock_module_0.puc_noscan_n ),
    .Y(_00108_)
  );
  AOI21X1 _05777_ (
    .A( clock_module_0.dbg_rst ),
    .B(_00108_),
    .C( clock_module_0.dbg_cpu_reset ),
    .Y( clock_module_0.sync_cell_puc.data_in )
  );
  NOR2X1 _05778_ (
    .A(_05632_),
    .B(1'h0),
    .Y(_00109_)
  );
  NAND3X1 _05779_ (
    .A(_00100_),
    .B(_05659_),
    .C(_00109_),
    .Y(_00110_)
  );
  INVX1 _05780_ (
    .A(_00110_),
    .Y(_00111_)
  );
  NOR2X1 _05781_ (
    .A(_05641_),
    .B(_05640_),
    .Y(_00112_)
  );
  NOR2X1 _05782_ (
    .A(_05631_),
    .B(_05642_),
    .Y(_00113_)
  );
  NAND2X1 _05783_ (
    .A(_00112_),
    .B(_00113_),
    .Y(_00114_)
  );
  NAND2X1 _05784_ (
    .A(_00098_),
    .B(_05636_),
    .Y(_00115_)
  );
  NAND2X1 _05785_ (
    .A(_00099_),
    .B(_05638_),
    .Y(_00116_)
  );
  NOR3X1 _05786_ (
    .A(_00114_),
    .B(_00115_),
    .C(_00116_),
    .Y(_00117_)
  );
  NOR2X1 _05787_ (
    .A(_05661_),
    .B(_05660_),
    .Y(_00118_)
  );
  NAND3X1 _05788_ (
    .A(_00111_),
    .B(_00117_),
    .C(_00118_),
    .Y(_00119_)
  );
  NOR2X1 _05789_ (
    .A(_05634_),
    .B(_05630_),
    .Y(_00120_)
  );
  AND2X1 _05790_ (
    .A(_05635_),
    .B(_00120_),
    .Y(_00121_)
  );
  NAND2X1 _05791_ (
    .A(_05635_),
    .B(_00120_),
    .Y(_00062_)
  );
  NOR2X1 _05792_ (
    .A(_00119_),
    .B(_00062_),
    .Y(_00063_)
  );
  AND2X1 _05793_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B(_00063_),
    .Y( clock_module_0.bcsctl2_rd_1_ )
  );
  AND2X1 _05794_ (
    .A( clock_module_0.bcsctl2_2_ ),
    .B(_00063_),
    .Y( clock_module_0.bcsctl2_rd_2_ )
  );
  AND2X1 _05795_ (
    .A( clock_module_0.bcsctl2_3_ ),
    .B(_00063_),
    .Y( clock_module_0.bcsctl2_rd_3_ )
  );
  NAND2X1 _05796_ (
    .A(_05634_),
    .B(_05630_),
    .Y(_00064_)
  );
  NOR2X1 _05797_ (
    .A(_05635_),
    .B(_00064_),
    .Y(_00065_)
  );
  NOR3X1 _05798_ (
    .A(_05635_),
    .B(_00119_),
    .C(_00064_),
    .Y(_00066_)
  );
  AND2X1 _05799_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B(_00066_),
    .Y( clock_module_0.bcsctl1_rd_12_ )
  );
  AND2X1 _05800_ (
    .A( clock_module_0.bcsctl1_5_ ),
    .B(_00066_),
    .Y( clock_module_0.bcsctl1_rd_13_ )
  );
  OAI21X1 _05801_ (
    .A(_00102_),
    .B( clock_module_0.aclk_div_2_ ),
    .C( clock_module_0.aclk_div_1_ ),
    .Y(_00067_)
  );
  OR2X1 _05802_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B( clock_module_0.bcsctl1_5_ ),
    .Y(_00068_)
  );
  OAI21X1 _05803_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B( clock_module_0.bcsctl1_5_ ),
    .C(_00097_),
    .Y(_00069_)
  );
  NAND2X1 _05804_ (
    .A(_00103_),
    .B( clock_module_0.lfxt_clk_s ),
    .Y(_00070_)
  );
  NOR2X1 _05805_ (
    .A( clock_module_0.oscoff ),
    .B(_00070_),
    .Y(_00071_)
  );
  NAND3X1 _05806_ (
    .A(_00103_),
    .B( clock_module_0.lfxt_clk_s ),
    .C(_00104_),
    .Y(_00072_)
  );
  NAND3X1 _05807_ (
    .A(cpu_en),
    .B(_00069_),
    .C(_00071_),
    .Y(_00073_)
  );
  AOI21X1 _05808_ (
    .A( clock_module_0.bcsctl1_5_ ),
    .B(_00067_),
    .C(_00073_),
    .Y(_00048_)
  );
  AOI21X1 _05809_ (
    .A( clock_module_0.bcsctl2_3_ ),
    .B(_00072_),
    .C( clock_module_0.scg1 ),
    .Y(_00074_)
  );
  AOI21X1 _05810_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B(_00107_),
    .C(_00106_),
    .Y(_00075_)
  );
  OR2X1 _05811_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B( clock_module_0.bcsctl2_2_ ),
    .Y(_00076_)
  );
  OAI21X1 _05812_ (
    .A(_00101_),
    .B(_00075_),
    .C( clock_module_0.smclk_div_0_ ),
    .Y(_00077_)
  );
  NAND2X1 _05813_ (
    .A(cpu_en),
    .B(_00074_),
    .Y(_00078_)
  );
  AOI21X1 _05814_ (
    .A(_00076_),
    .B(_00077_),
    .C(_00078_),
    .Y(_00049_)
  );
  OR2X1 _05815_ (
    .A( clock_module_0.wdt_reset ),
    .B( clock_module_0.por ),
    .Y( clock_module_0.puc_a )
  );
  NOR2X1 _05816_ (
    .A(_05641_),
    .B(_05642_),
    .Y(_00079_)
  );
  NAND3X1 _05817_ (
    .A(_00098_),
    .B(_00099_),
    .C(_00079_),
    .Y(_00080_)
  );
  NOR2X1 _05818_ (
    .A(_05640_),
    .B(_05631_),
    .Y(_00081_)
  );
  NAND3X1 _05819_ (
    .A(_05636_),
    .B(_05638_),
    .C(_00081_),
    .Y(_00082_)
  );
  NOR3X1 _05820_ (
    .A(_00110_),
    .B(_00080_),
    .C(_00082_),
    .Y(_00083_)
  );
  NAND3X1 _05821_ (
    .A(_05660_),
    .B(_00121_),
    .C(_00083_),
    .Y(_00084_)
  );
  MUX2X1 _05822_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B(_05650_),
    .S(_00084_),
    .Y(_00085_)
  );
  INVX1 _05823_ (
    .A(_00085_),
    .Y(_00051_)
  );
  MUX2X1 _05824_ (
    .A( clock_module_0.bcsctl2_2_ ),
    .B(_05651_),
    .S(_00084_),
    .Y(_00086_)
  );
  INVX1 _05825_ (
    .A(_00086_),
    .Y(_00052_)
  );
  MUX2X1 _05826_ (
    .A( clock_module_0.bcsctl2_3_ ),
    .B(_05652_),
    .S(_00084_),
    .Y(_00087_)
  );
  INVX1 _05827_ (
    .A(_00087_),
    .Y(_00053_)
  );
  OAI21X1 _05828_ (
    .A( clock_module_0.bcsctl2_1_ ),
    .B( clock_module_0.bcsctl2_2_ ),
    .C(_00074_),
    .Y(_00088_)
  );
  NAND3X1 _05829_ (
    .A( clock_module_0.smclk_div_0_ ),
    .B(_00074_),
    .C(_00076_),
    .Y(_00089_)
  );
  XNOR2X1 _05830_ (
    .A( clock_module_0.smclk_div_0_ ),
    .B(_00088_),
    .Y(_00054_)
  );
  NOR2X1 _05831_ (
    .A(_00106_),
    .B(_00089_),
    .Y(_00090_)
  );
  XNOR2X1 _05832_ (
    .A( clock_module_0.smclk_div_1_ ),
    .B(_00089_),
    .Y(_00055_)
  );
  XNOR2X1 _05833_ (
    .A(_00107_),
    .B(_00090_),
    .Y(_00056_)
  );
  OAI21X1 _05834_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B( clock_module_0.bcsctl1_5_ ),
    .C(_00071_),
    .Y(_00091_)
  );
  NAND3X1 _05835_ (
    .A( clock_module_0.aclk_div_0_ ),
    .B(_00068_),
    .C(_00071_),
    .Y(_00092_)
  );
  XNOR2X1 _05836_ (
    .A( clock_module_0.aclk_div_0_ ),
    .B(_00091_),
    .Y(_00057_)
  );
  NOR2X1 _05837_ (
    .A(_00105_),
    .B(_00092_),
    .Y(_00093_)
  );
  XNOR2X1 _05838_ (
    .A( clock_module_0.aclk_div_1_ ),
    .B(_00092_),
    .Y(_00058_)
  );
  XOR2X1 _05839_ (
    .A( clock_module_0.aclk_div_2_ ),
    .B(_00093_),
    .Y(_00059_)
  );
  NAND3X1 _05840_ (
    .A(_05661_),
    .B(_00065_),
    .C(_00083_),
    .Y(_00094_)
  );
  MUX2X1 _05841_ (
    .A( clock_module_0.bcsctl1_4_ ),
    .B(_05646_),
    .S(_00094_),
    .Y(_00095_)
  );
  INVX1 _05842_ (
    .A(_00095_),
    .Y(_00060_)
  );
  MUX2X1 _05843_ (
    .A( clock_module_0.bcsctl1_5_ ),
    .B(_05647_),
    .S(_00094_),
    .Y(_00096_)
  );
  INVX1 _05844_ (
    .A(_00096_),
    .Y(_00061_)
  );
  DFFSR _05845_ (
    .CLK(dco_clk),
    .D( clock_module_0.dbg_rst_nxt ),
    .Q( clock_module_0.dbg_rst ),
    .R(1'h1),
    .S(_00050_)
  );
  DFFSR _05846_ (
    .CLK(dco_clk),
    .D(_00051_),
    .Q( clock_module_0.bcsctl2_1_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05847_ (
    .CLK(dco_clk),
    .D(_00052_),
    .Q( clock_module_0.bcsctl2_2_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05848_ (
    .CLK(dco_clk),
    .D(_00053_),
    .Q( clock_module_0.bcsctl2_3_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05849_ (
    .CLK(dco_clk),
    .D(_00049_),
    .Q(_05696_),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05850_ (
    .CLK(dco_clk),
    .D(_00048_),
    .Q(_05581_),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05851_ (
    .CLK(dco_clk),
    .D(_00054_),
    .Q( clock_module_0.smclk_div_0_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05852_ (
    .CLK(dco_clk),
    .D(_00055_),
    .Q( clock_module_0.smclk_div_1_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05853_ (
    .CLK(dco_clk),
    .D(_00056_),
    .Q( clock_module_0.smclk_div_2_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05854_ (
    .CLK(dco_clk),
    .D( clock_module_0.lfxt_clk_s ),
    .Q( clock_module_0.lfxt_clk_dly ),
    .R(_00050_),
    .S(1'h1)
  );
  DFFSR _05855_ (
    .CLK(dco_clk),
    .D(_00057_),
    .Q( clock_module_0.aclk_div_0_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05856_ (
    .CLK(dco_clk),
    .D(_00058_),
    .Q( clock_module_0.aclk_div_1_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05857_ (
    .CLK(dco_clk),
    .D(_00059_),
    .Q( clock_module_0.aclk_div_2_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05858_ (
    .CLK(dco_clk),
    .D(_00060_),
    .Q( clock_module_0.bcsctl1_4_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _05859_ (
    .CLK(dco_clk),
    .D(_00061_),
    .Q( clock_module_0.bcsctl1_5_ ),
    .R( clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  INVX1 _05860_ (
    .A( clock_module_0.por ),
    .Y(_00122_)
  );
  DFFSR _05861_ (
    .CLK(dco_clk),
    .D(lfxt_clk),
    .Q( clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .R(_00122_),
    .S(1'h1)
  );
  DFFSR _05862_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .Q( clock_module_0.lfxt_clk_s ),
    .R(_00122_),
    .S(1'h1)
  );
  INVX1 _05863_ (
    .A( clock_module_0.puc_a ),
    .Y(_00123_)
  );
  DFFSR _05864_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_cell_puc.data_in ),
    .Q( clock_module_0.sync_cell_puc.data_sync_0_ ),
    .R(_00123_),
    .S(1'h1)
  );
  DFFSR _05865_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_cell_puc.data_sync_0_ ),
    .Q( clock_module_0.puc_noscan_n ),
    .R(_00123_),
    .S(1'h1)
  );
  INVX1 _05866_ (
    .A( clock_module_0.por_a ),
    .Y(_00124_)
  );
  DFFSR _05867_ (
    .CLK(dco_clk),
    .D(1'h0),
    .Q( clock_module_0.sync_reset_por.data_sync_0_ ),
    .R(1'h1),
    .S(_00124_)
  );
  DFFSR _05868_ (
    .CLK(dco_clk),
    .D( clock_module_0.sync_reset_por.data_sync_0_ ),
    .Q( clock_module_0.por ),
    .R(1'h1),
    .S(_00124_)
  );
  INVX1 _05869_ (
    .A( dbg_0.mem_cnt_8_ ),
    .Y(_00189_)
  );
  INVX1 _05870_ (
    .A( dbg_0.mem_cnt_13_ ),
    .Y(_00190_)
  );
  INVX1 _05871_ (
    .A( dbg_0.mem_cnt_12_ ),
    .Y(_00191_)
  );
  INVX1 _05872_ (
    .A( dbg_0.mem_cnt_14_ ),
    .Y(_00192_)
  );
  INVX1 _05873_ (
    .A( dbg_0.mem_state_1_ ),
    .Y(_00193_)
  );
  INVX1 _05874_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_00194_)
  );
  INVX1 _05875_ (
    .A( dbg_0.dbg_addr_0_ ),
    .Y(_00195_)
  );
  INVX1 _05876_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00196_)
  );
  INVX1 _05877_ (
    .A( dbg_0.mem_ctl_1_ ),
    .Y(_00197_)
  );
  INVX1 _05878_ (
    .A( dbg_0.dbg_mem_rd_dly ),
    .Y(_00198_)
  );
  INVX1 _05879_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .Y(_00199_)
  );
  INVX1 _05880_ (
    .A( dbg_0.dbg_din_0_ ),
    .Y(_00200_)
  );
  INVX1 _05881_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .Y(_00201_)
  );
  INVX1 _05882_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .Y(_00202_)
  );
  INVX1 _05883_ (
    .A( dbg_0.dbg_mem_addr_4_ ),
    .Y(_00203_)
  );
  INVX1 _05884_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .Y(_00204_)
  );
  INVX1 _05885_ (
    .A( dbg_0.dbg_din_5_ ),
    .Y(_00205_)
  );
  INVX1 _05886_ (
    .A( dbg_0.dbg_din_7_ ),
    .Y(_00206_)
  );
  INVX1 _05887_ (
    .A( dbg_0.dbg_mem_addr_8_ ),
    .Y(_00207_)
  );
  INVX1 _05888_ (
    .A( dbg_0.dbg_din_8_ ),
    .Y(_00208_)
  );
  INVX1 _05889_ (
    .A( dbg_0.dbg_mem_addr_9_ ),
    .Y(_00209_)
  );
  INVX1 _05890_ (
    .A( dbg_0.dbg_din_9_ ),
    .Y(_00210_)
  );
  INVX1 _05891_ (
    .A( dbg_0.dbg_mem_addr_12_ ),
    .Y(_00211_)
  );
  INVX1 _05892_ (
    .A( dbg_0.dbg_din_13_ ),
    .Y(_00212_)
  );
  INVX1 _05893_ (
    .A( dbg_0.dbg_din_15_ ),
    .Y(_00213_)
  );
  INVX1 _05894_ (
    .A( dbg_0.mem_data_0_ ),
    .Y(_00214_)
  );
  INVX1 _05895_ (
    .A( dbg_0.mem_data_1_ ),
    .Y(_00215_)
  );
  INVX1 _05896_ (
    .A( dbg_0.mem_data_2_ ),
    .Y(_00216_)
  );
  INVX1 _05897_ (
    .A( dbg_0.mem_data_3_ ),
    .Y(_00217_)
  );
  INVX1 _05898_ (
    .A( dbg_0.mem_data_4_ ),
    .Y(_00218_)
  );
  INVX1 _05899_ (
    .A( dbg_0.mem_data_5_ ),
    .Y(_00219_)
  );
  INVX1 _05900_ (
    .A( dbg_0.mem_data_6_ ),
    .Y(_00220_)
  );
  INVX1 _05901_ (
    .A( dbg_0.mem_data_7_ ),
    .Y(_00221_)
  );
  INVX1 _05902_ (
    .A( dbg_0.mem_data_8_ ),
    .Y(_00222_)
  );
  INVX1 _05903_ (
    .A( dbg_0.mem_data_9_ ),
    .Y(_00223_)
  );
  INVX1 _05904_ (
    .A( dbg_0.mem_data_10_ ),
    .Y(_00224_)
  );
  INVX1 _05905_ (
    .A( dbg_0.mem_data_11_ ),
    .Y(_00225_)
  );
  INVX1 _05906_ (
    .A( dbg_0.mem_data_12_ ),
    .Y(_00226_)
  );
  INVX1 _05907_ (
    .A( dbg_0.mem_data_13_ ),
    .Y(_00227_)
  );
  INVX1 _05908_ (
    .A( dbg_0.mem_data_14_ ),
    .Y(_00228_)
  );
  INVX1 _05909_ (
    .A( dbg_0.mem_data_15_ ),
    .Y(_00229_)
  );
  INVX1 _05910_ (
    .A(cpu_en),
    .Y(_00230_)
  );
  INVX1 _05911_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00163_)
  );
  NOR2X1 _05912_ (
    .A( dbg_0.mem_cnt_5_ ),
    .B( dbg_0.mem_cnt_4_ ),
    .Y(_00231_)
  );
  OR2X1 _05913_ (
    .A( dbg_0.mem_cnt_5_ ),
    .B( dbg_0.mem_cnt_4_ ),
    .Y(_00232_)
  );
  NOR2X1 _05914_ (
    .A( dbg_0.mem_cnt_7_ ),
    .B( dbg_0.mem_cnt_6_ ),
    .Y(_00233_)
  );
  OR2X1 _05915_ (
    .A( dbg_0.mem_cnt_6_ ),
    .B(_00232_),
    .Y(_00234_)
  );
  NAND2X1 _05916_ (
    .A(_00231_),
    .B(_00233_),
    .Y(_00235_)
  );
  NOR2X1 _05917_ (
    .A( dbg_0.mem_cnt_0_ ),
    .B( dbg_0.mem_cnt_3_ ),
    .Y(_00236_)
  );
  NOR2X1 _05918_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B( dbg_0.mem_cnt_2_ ),
    .Y(_00237_)
  );
  OR2X1 _05919_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B( dbg_0.mem_cnt_2_ ),
    .Y(_00238_)
  );
  NAND2X1 _05920_ (
    .A(_00236_),
    .B(_00237_),
    .Y(_00239_)
  );
  NOR2X1 _05921_ (
    .A( dbg_0.mem_cnt_9_ ),
    .B( dbg_0.mem_cnt_8_ ),
    .Y(_00240_)
  );
  NOR2X1 _05922_ (
    .A( dbg_0.mem_cnt_11_ ),
    .B( dbg_0.mem_cnt_10_ ),
    .Y(_00241_)
  );
  NAND2X1 _05923_ (
    .A(_00240_),
    .B(_00241_),
    .Y(_00242_)
  );
  NOR2X1 _05924_ (
    .A( dbg_0.mem_cnt_15_ ),
    .B( dbg_0.mem_cnt_14_ ),
    .Y(_00243_)
  );
  NAND3X1 _05925_ (
    .A(_00236_),
    .B(_00240_),
    .C(_00241_),
    .Y(_00244_)
  );
  NAND3X1 _05926_ (
    .A(_00191_),
    .B(_00237_),
    .C(_00243_),
    .Y(_00245_)
  );
  NAND3X1 _05927_ (
    .A(_00190_),
    .B(_00231_),
    .C(_00233_),
    .Y(_00246_)
  );
  NOR3X1 _05928_ (
    .A(_00244_),
    .B(_00245_),
    .C(_00246_),
    .Y(_00247_)
  );
  INVX1 _05929_ (
    .A(_00247_),
    .Y(_00248_)
  );
  AOI21X1 _05930_ (
    .A( dbg_0.mem_start ),
    .B(_00247_),
    .C( dbg_0.mem_startb ),
    .Y(_00249_)
  );
  INVX1 _05931_ (
    .A(_00249_),
    .Y(_00250_)
  );
  NAND2X1 _05932_ (
    .A(_00193_),
    .B(_00250_),
    .Y(_00251_)
  );
  OAI21X1 _05933_ (
    .A( dbg_0.mem_state_0_ ),
    .B(_00250_),
    .C(_00193_),
    .Y(_00252_)
  );
  AOI21X1 _05934_ (
    .A( dbg_0.mem_state_0_ ),
    .B( dbg_0.cpu_stat_full_0_ ),
    .C(_00252_),
    .Y( dbg_0.mem_state_nxt_0_ )
  );
  AND2X1 _05935_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B( dbg_0.dbg_mem_addr_0_ ),
    .Y(_00253_)
  );
  NAND2X1 _05936_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B( dbg_0.dbg_mem_addr_0_ ),
    .Y(_00254_)
  );
  NOR2X1 _05937_ (
    .A(_00193_),
    .B( dbg_0.mem_ctl_2_ ),
    .Y( dbg_0.dbg_mem_en )
  );
  NOR2X1 _05938_ (
    .A(_00193_),
    .B(_00197_),
    .Y(_00255_)
  );
  NAND2X1 _05939_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B( dbg_0.dbg_mem_en ),
    .Y(_00256_)
  );
  NOR2X1 _05940_ (
    .A(_00253_),
    .B(_00256_),
    .Y( dbg_0.dbg_mem_wr_0_ )
  );
  AOI21X1 _05941_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00199_),
    .C(_00256_),
    .Y( dbg_0.dbg_mem_wr_1_ )
  );
  NOR2X1 _05942_ (
    .A(_00194_),
    .B(_00252_),
    .Y( dbg_0.mem_state_nxt_1_ )
  );
  OAI21X1 _05943_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B( dbg_0.dbg_rd_rdy ),
    .C(_00247_),
    .Y(_00257_)
  );
  INVX1 _05944_ (
    .A(_00257_),
    .Y( dbg_0.dbg_i2c_0.mem_burst_end )
  );
  AND2X1 _05945_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B(_00255_),
    .Y( dbg_0.dbg_reg_wr )
  );
  NOR2X1 _05946_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_addr_1_ ),
    .Y(_00258_)
  );
  NAND2X1 _05947_ (
    .A( dbg_0.dbg_addr_0_ ),
    .B(_00258_),
    .Y(_00259_)
  );
  OR2X1 _05948_ (
    .A( dbg_0.dbg_addr_4_ ),
    .B( dbg_0.dbg_addr_5_ ),
    .Y(_00260_)
  );
  NOR2X1 _05949_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_addr_2_ ),
    .Y(_00261_)
  );
  OAI21X1 _05950_ (
    .A( dbg_0.dbg_addr_3_ ),
    .B(_00260_),
    .C(_00196_),
    .Y(_00262_)
  );
  OAI21X1 _05951_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_addr_2_ ),
    .C(_00262_),
    .Y(_00263_)
  );
  NOR2X1 _05952_ (
    .A(_00259_),
    .B(_00263_),
    .Y(_00264_)
  );
  AND2X1 _05953_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00264_),
    .Y(_00265_)
  );
  NAND2X1 _05954_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00264_),
    .Y(_00266_)
  );
  NOR2X1 _05955_ (
    .A( dbg_0.dbg_rd_rdy ),
    .B(_00255_),
    .Y(_00267_)
  );
  NOR2X1 _05956_ (
    .A(_00196_),
    .B(_00267_),
    .Y(_00268_)
  );
  OAI21X1 _05957_ (
    .A( dbg_0.dbg_rd_rdy ),
    .B(_00255_),
    .C( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00269_)
  );
  NOR2X1 _05958_ (
    .A(_00247_),
    .B(_00269_),
    .Y(_00270_)
  );
  NAND2X1 _05959_ (
    .A(_00248_),
    .B(_00268_),
    .Y(_00271_)
  );
  NOR2X1 _05960_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B( dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00272_)
  );
  OR2X1 _05961_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B( dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00273_)
  );
  NAND3X1 _05962_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .B(_00270_),
    .C(_00273_),
    .Y(_00274_)
  );
  OAI21X1 _05963_ (
    .A(_00271_),
    .B(_00272_),
    .C(_00199_),
    .Y(_00275_)
  );
  NAND2X1 _05964_ (
    .A(_00274_),
    .B(_00275_),
    .Y(_00276_)
  );
  NAND2X1 _05965_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00265_),
    .Y(_00277_)
  );
  OAI21X1 _05966_ (
    .A(_00265_),
    .B(_00276_),
    .C(_00277_),
    .Y(_00129_)
  );
  NOR3X1 _05967_ (
    .A(_00247_),
    .B(_00269_),
    .C(_00273_),
    .Y(_00278_)
  );
  NAND2X1 _05968_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .B(_00278_),
    .Y(_00279_)
  );
  XNOR2X1 _05969_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .B(_00278_),
    .Y(_00280_)
  );
  XNOR2X1 _05970_ (
    .A(_00274_),
    .B(_00280_),
    .Y(_00281_)
  );
  NAND2X1 _05971_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00265_),
    .Y(_00282_)
  );
  OAI21X1 _05972_ (
    .A(_00265_),
    .B(_00281_),
    .C(_00282_),
    .Y(_00136_)
  );
  OAI21X1 _05973_ (
    .A(_00274_),
    .B(_00280_),
    .C(_00279_),
    .Y(_00283_)
  );
  AND2X1 _05974_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00283_),
    .Y(_00284_)
  );
  NAND2X1 _05975_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00283_),
    .Y(_00285_)
  );
  OAI21X1 _05976_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00283_),
    .C(_00266_),
    .Y(_00286_)
  );
  NAND2X1 _05977_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00265_),
    .Y(_00287_)
  );
  OAI21X1 _05978_ (
    .A(_00284_),
    .B(_00286_),
    .C(_00287_),
    .Y(_00137_)
  );
  NAND3X1 _05979_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B( dbg_0.dbg_mem_addr_3_ ),
    .C(_00283_),
    .Y(_00288_)
  );
  XOR2X1 _05980_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_00285_),
    .Y(_00289_)
  );
  NAND2X1 _05981_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00265_),
    .Y(_00290_)
  );
  OAI21X1 _05982_ (
    .A(_00265_),
    .B(_00289_),
    .C(_00290_),
    .Y(_00138_)
  );
  NAND2X1 _05983_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00265_),
    .Y(_00291_)
  );
  NOR2X1 _05984_ (
    .A(_00203_),
    .B(_00288_),
    .Y(_00292_)
  );
  XNOR2X1 _05985_ (
    .A(_00203_),
    .B(_00288_),
    .Y(_00293_)
  );
  OAI21X1 _05986_ (
    .A(_00265_),
    .B(_00293_),
    .C(_00291_),
    .Y(_00139_)
  );
  NOR2X1 _05987_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .B(_00292_),
    .Y(_00294_)
  );
  NOR3X1 _05988_ (
    .A(_00203_),
    .B(_00204_),
    .C(_00288_),
    .Y(_00295_)
  );
  OR2X1 _05989_ (
    .A(_00265_),
    .B(_00295_),
    .Y(_00296_)
  );
  OAI22X1 _05990_ (
    .A(_00205_),
    .B(_00266_),
    .C(_00294_),
    .D(_00296_),
    .Y(_00140_)
  );
  NAND2X1 _05991_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00265_),
    .Y(_00297_)
  );
  AND2X1 _05992_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00295_),
    .Y(_00298_)
  );
  OAI21X1 _05993_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00295_),
    .C(_00266_),
    .Y(_00299_)
  );
  OAI21X1 _05994_ (
    .A(_00298_),
    .B(_00299_),
    .C(_00297_),
    .Y(_00141_)
  );
  NAND3X1 _05995_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B( dbg_0.dbg_mem_addr_7_ ),
    .C(_00295_),
    .Y(_00300_)
  );
  AOI21X1 _05996_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00295_),
    .C( dbg_0.dbg_mem_addr_7_ ),
    .Y(_00301_)
  );
  NOR2X1 _05997_ (
    .A(_00265_),
    .B(_00301_),
    .Y(_00302_)
  );
  NAND2X1 _05998_ (
    .A(_00300_),
    .B(_00302_),
    .Y(_00303_)
  );
  OAI21X1 _05999_ (
    .A(_00206_),
    .B(_00266_),
    .C(_00303_),
    .Y(_00142_)
  );
  NAND2X1 _06000_ (
    .A( dbg_0.dbg_din_8_ ),
    .B(_00265_),
    .Y(_00304_)
  );
  XNOR2X1 _06001_ (
    .A(_00207_),
    .B(_00300_),
    .Y(_00305_)
  );
  OAI21X1 _06002_ (
    .A(_00265_),
    .B(_00305_),
    .C(_00304_),
    .Y(_00143_)
  );
  OAI21X1 _06003_ (
    .A(_00207_),
    .B(_00300_),
    .C(_00209_),
    .Y(_00306_)
  );
  NOR3X1 _06004_ (
    .A(_00207_),
    .B(_00209_),
    .C(_00300_),
    .Y(_00307_)
  );
  NOR2X1 _06005_ (
    .A(_00265_),
    .B(_00307_),
    .Y(_00308_)
  );
  NAND2X1 _06006_ (
    .A(_00306_),
    .B(_00308_),
    .Y(_00309_)
  );
  OAI21X1 _06007_ (
    .A(_00210_),
    .B(_00266_),
    .C(_00309_),
    .Y(_00144_)
  );
  NAND2X1 _06008_ (
    .A( dbg_0.dbg_din_10_ ),
    .B(_00265_),
    .Y(_00310_)
  );
  NAND2X1 _06009_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B(_00307_),
    .Y(_00311_)
  );
  XNOR2X1 _06010_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B(_00307_),
    .Y(_00312_)
  );
  OAI21X1 _06011_ (
    .A(_00265_),
    .B(_00312_),
    .C(_00310_),
    .Y(_00130_)
  );
  NAND2X1 _06012_ (
    .A( dbg_0.dbg_din_11_ ),
    .B(_00265_),
    .Y(_00313_)
  );
  NAND3X1 _06013_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B( dbg_0.dbg_mem_addr_11_ ),
    .C(_00307_),
    .Y(_00314_)
  );
  XOR2X1 _06014_ (
    .A( dbg_0.dbg_mem_addr_11_ ),
    .B(_00311_),
    .Y(_00315_)
  );
  OAI21X1 _06015_ (
    .A(_00265_),
    .B(_00315_),
    .C(_00313_),
    .Y(_00131_)
  );
  NAND2X1 _06016_ (
    .A( dbg_0.dbg_din_12_ ),
    .B(_00265_),
    .Y(_00316_)
  );
  NOR2X1 _06017_ (
    .A(_00211_),
    .B(_00314_),
    .Y(_00317_)
  );
  XNOR2X1 _06018_ (
    .A(_00211_),
    .B(_00314_),
    .Y(_00318_)
  );
  OAI21X1 _06019_ (
    .A(_00265_),
    .B(_00318_),
    .C(_00316_),
    .Y(_00132_)
  );
  NAND2X1 _06020_ (
    .A( dbg_0.dbg_din_13_ ),
    .B(_00265_),
    .Y(_00319_)
  );
  NAND2X1 _06021_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B(_00317_),
    .Y(_00320_)
  );
  XNOR2X1 _06022_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B(_00317_),
    .Y(_00321_)
  );
  OAI21X1 _06023_ (
    .A(_00265_),
    .B(_00321_),
    .C(_00319_),
    .Y(_00133_)
  );
  NAND2X1 _06024_ (
    .A( dbg_0.dbg_din_14_ ),
    .B(_00265_),
    .Y(_00322_)
  );
  NAND3X1 _06025_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B( dbg_0.dbg_mem_addr_14_ ),
    .C(_00317_),
    .Y(_00323_)
  );
  XOR2X1 _06026_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .B(_00320_),
    .Y(_00324_)
  );
  OAI21X1 _06027_ (
    .A(_00265_),
    .B(_00324_),
    .C(_00322_),
    .Y(_00134_)
  );
  XOR2X1 _06028_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .B(_00323_),
    .Y(_00325_)
  );
  MUX2X1 _06029_ (
    .A(_00213_),
    .B(_00325_),
    .S(_00265_),
    .Y(_00135_)
  );
  NAND3X1 _06030_ (
    .A( dbg_0.dbg_addr_0_ ),
    .B(_00196_),
    .C( dbg_0.dbg_addr_1_ ),
    .Y(_00326_)
  );
  NOR2X1 _06031_ (
    .A(_00263_),
    .B(_00326_),
    .Y(_00327_)
  );
  AND2X1 _06032_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00327_),
    .Y(_00328_)
  );
  NAND2X1 _06033_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00327_),
    .Y(_00329_)
  );
  OR2X1 _06034_ (
    .A( dbg_0.mem_cnt_0_ ),
    .B(_00271_),
    .Y(_00330_)
  );
  OAI21X1 _06035_ (
    .A(_00247_),
    .B(_00269_),
    .C( dbg_0.mem_cnt_0_ ),
    .Y(_00331_)
  );
  AND2X1 _06036_ (
    .A(_00330_),
    .B(_00331_),
    .Y(_00332_)
  );
  NAND2X1 _06037_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00328_),
    .Y(_00333_)
  );
  OAI21X1 _06038_ (
    .A(_00328_),
    .B(_00332_),
    .C(_00333_),
    .Y(_00145_)
  );
  NOR2X1 _06039_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B(_00330_),
    .Y(_00334_)
  );
  XOR2X1 _06040_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B(_00330_),
    .Y(_00335_)
  );
  NAND2X1 _06041_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00328_),
    .Y(_00336_)
  );
  OAI21X1 _06042_ (
    .A(_00328_),
    .B(_00335_),
    .C(_00336_),
    .Y(_00152_)
  );
  XNOR2X1 _06043_ (
    .A( dbg_0.mem_cnt_2_ ),
    .B(_00334_),
    .Y(_00337_)
  );
  NAND2X1 _06044_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00328_),
    .Y(_00338_)
  );
  OAI21X1 _06045_ (
    .A(_00328_),
    .B(_00337_),
    .C(_00338_),
    .Y(_00153_)
  );
  OR2X1 _06046_ (
    .A(_00239_),
    .B(_00271_),
    .Y(_00339_)
  );
  OAI21X1 _06047_ (
    .A(_00238_),
    .B(_00330_),
    .C( dbg_0.mem_cnt_3_ ),
    .Y(_00340_)
  );
  AND2X1 _06048_ (
    .A(_00339_),
    .B(_00340_),
    .Y(_00341_)
  );
  NAND2X1 _06049_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00328_),
    .Y(_00342_)
  );
  OAI21X1 _06050_ (
    .A(_00328_),
    .B(_00341_),
    .C(_00342_),
    .Y(_00154_)
  );
  XOR2X1 _06051_ (
    .A( dbg_0.mem_cnt_4_ ),
    .B(_00339_),
    .Y(_00343_)
  );
  NAND2X1 _06052_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00328_),
    .Y(_00344_)
  );
  OAI21X1 _06053_ (
    .A(_00328_),
    .B(_00343_),
    .C(_00344_),
    .Y(_00155_)
  );
  OAI21X1 _06054_ (
    .A( dbg_0.mem_cnt_4_ ),
    .B(_00339_),
    .C( dbg_0.mem_cnt_5_ ),
    .Y(_00345_)
  );
  OAI21X1 _06055_ (
    .A(_00232_),
    .B(_00339_),
    .C(_00345_),
    .Y(_00346_)
  );
  NAND2X1 _06056_ (
    .A(_00329_),
    .B(_00346_),
    .Y(_00347_)
  );
  OAI21X1 _06057_ (
    .A(_00205_),
    .B(_00329_),
    .C(_00347_),
    .Y(_00156_)
  );
  OR2X1 _06058_ (
    .A(_00234_),
    .B(_00339_),
    .Y(_00348_)
  );
  OAI21X1 _06059_ (
    .A(_00232_),
    .B(_00339_),
    .C( dbg_0.mem_cnt_6_ ),
    .Y(_00349_)
  );
  AND2X1 _06060_ (
    .A(_00348_),
    .B(_00349_),
    .Y(_00350_)
  );
  NAND2X1 _06061_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00328_),
    .Y(_00351_)
  );
  OAI21X1 _06062_ (
    .A(_00328_),
    .B(_00350_),
    .C(_00351_),
    .Y(_00157_)
  );
  NOR2X1 _06063_ (
    .A( dbg_0.dbg_din_7_ ),
    .B(_00329_),
    .Y(_00352_)
  );
  XOR2X1 _06064_ (
    .A( dbg_0.mem_cnt_7_ ),
    .B(_00348_),
    .Y(_00353_)
  );
  AOI21X1 _06065_ (
    .A(_00329_),
    .B(_00353_),
    .C(_00352_),
    .Y(_00158_)
  );
  OAI21X1 _06066_ (
    .A(_00235_),
    .B(_00239_),
    .C(_00268_),
    .Y(_00354_)
  );
  NAND2X1 _06067_ (
    .A(_00270_),
    .B(_00354_),
    .Y(_00355_)
  );
  OR2X1 _06068_ (
    .A( dbg_0.mem_cnt_8_ ),
    .B(_00354_),
    .Y(_00356_)
  );
  XNOR2X1 _06069_ (
    .A(_00189_),
    .B(_00355_),
    .Y(_00357_)
  );
  MUX2X1 _06070_ (
    .A(_00208_),
    .B(_00357_),
    .S(_00328_),
    .Y(_00159_)
  );
  OAI21X1 _06071_ (
    .A(_00189_),
    .B(_00271_),
    .C(_00356_),
    .Y(_00358_)
  );
  XNOR2X1 _06072_ (
    .A( dbg_0.mem_cnt_9_ ),
    .B(_00270_),
    .Y(_00359_)
  );
  XOR2X1 _06073_ (
    .A(_00358_),
    .B(_00359_),
    .Y(_00360_)
  );
  MUX2X1 _06074_ (
    .A(_00210_),
    .B(_00360_),
    .S(_00328_),
    .Y(_00160_)
  );
  OR2X1 _06075_ (
    .A(_00356_),
    .B(_00359_),
    .Y(_00361_)
  );
  OAI21X1 _06076_ (
    .A( dbg_0.mem_cnt_9_ ),
    .B( dbg_0.mem_cnt_8_ ),
    .C(_00270_),
    .Y(_00362_)
  );
  OAI21X1 _06077_ (
    .A(_00356_),
    .B(_00359_),
    .C(_00362_),
    .Y(_00363_)
  );
  XNOR2X1 _06078_ (
    .A( dbg_0.mem_cnt_10_ ),
    .B(_00270_),
    .Y(_00364_)
  );
  AOI21X1 _06079_ (
    .A(_00361_),
    .B(_00362_),
    .C(_00364_),
    .Y(_00365_)
  );
  XOR2X1 _06080_ (
    .A(_00363_),
    .B(_00364_),
    .Y(_00366_)
  );
  NAND2X1 _06081_ (
    .A( dbg_0.dbg_din_10_ ),
    .B(_00328_),
    .Y(_00367_)
  );
  OAI21X1 _06082_ (
    .A(_00328_),
    .B(_00366_),
    .C(_00367_),
    .Y(_00146_)
  );
  NOR2X1 _06083_ (
    .A( dbg_0.dbg_din_11_ ),
    .B(_00329_),
    .Y(_00368_)
  );
  AOI21X1 _06084_ (
    .A( dbg_0.mem_cnt_10_ ),
    .B(_00270_),
    .C(_00365_),
    .Y(_00369_)
  );
  XNOR2X1 _06085_ (
    .A( dbg_0.mem_cnt_11_ ),
    .B(_00270_),
    .Y(_00370_)
  );
  XNOR2X1 _06086_ (
    .A(_00369_),
    .B(_00370_),
    .Y(_00371_)
  );
  AOI21X1 _06087_ (
    .A(_00329_),
    .B(_00371_),
    .C(_00368_),
    .Y(_00147_)
  );
  NAND2X1 _06088_ (
    .A( dbg_0.dbg_din_12_ ),
    .B(_00328_),
    .Y(_00372_)
  );
  NAND2X1 _06089_ (
    .A(_00242_),
    .B(_00268_),
    .Y(_00373_)
  );
  OR2X1 _06090_ (
    .A(_00364_),
    .B(_00370_),
    .Y(_00374_)
  );
  OAI21X1 _06091_ (
    .A(_00361_),
    .B(_00374_),
    .C(_00373_),
    .Y(_00375_)
  );
  XNOR2X1 _06092_ (
    .A(_00191_),
    .B(_00270_),
    .Y(_00376_)
  );
  XNOR2X1 _06093_ (
    .A(_00375_),
    .B(_00376_),
    .Y(_00377_)
  );
  OAI21X1 _06094_ (
    .A(_00328_),
    .B(_00377_),
    .C(_00372_),
    .Y(_00148_)
  );
  AOI22X1 _06095_ (
    .A( dbg_0.mem_cnt_12_ ),
    .B(_00268_),
    .C(_00375_),
    .D(_00376_),
    .Y(_00378_)
  );
  OAI21X1 _06096_ (
    .A(_00247_),
    .B(_00269_),
    .C(_00190_),
    .Y(_00379_)
  );
  OAI21X1 _06097_ (
    .A(_00190_),
    .B(_00269_),
    .C(_00379_),
    .Y(_00380_)
  );
  AOI21X1 _06098_ (
    .A(_00378_),
    .B(_00380_),
    .C(_00328_),
    .Y(_00381_)
  );
  OAI21X1 _06099_ (
    .A(_00378_),
    .B(_00380_),
    .C(_00381_),
    .Y(_00382_)
  );
  OAI21X1 _06100_ (
    .A(_00212_),
    .B(_00329_),
    .C(_00382_),
    .Y(_00149_)
  );
  NAND2X1 _06101_ (
    .A( dbg_0.dbg_din_14_ ),
    .B(_00328_),
    .Y(_00383_)
  );
  XNOR2X1 _06102_ (
    .A(_00192_),
    .B(_00270_),
    .Y(_00384_)
  );
  OAI21X1 _06103_ (
    .A(_00190_),
    .B(_00271_),
    .C(_00378_),
    .Y(_00385_)
  );
  NAND2X1 _06104_ (
    .A(_00384_),
    .B(_00385_),
    .Y(_00386_)
  );
  XNOR2X1 _06105_ (
    .A(_00384_),
    .B(_00385_),
    .Y(_00387_)
  );
  OAI21X1 _06106_ (
    .A(_00328_),
    .B(_00387_),
    .C(_00383_),
    .Y(_00150_)
  );
  OAI21X1 _06107_ (
    .A(_00192_),
    .B(_00271_),
    .C(_00386_),
    .Y(_00388_)
  );
  XOR2X1 _06108_ (
    .A( dbg_0.mem_cnt_15_ ),
    .B(_00270_),
    .Y(_00389_)
  );
  XNOR2X1 _06109_ (
    .A(_00388_),
    .B(_00389_),
    .Y(_00390_)
  );
  NAND2X1 _06110_ (
    .A( dbg_0.dbg_din_15_ ),
    .B(_00328_),
    .Y(_00391_)
  );
  OAI21X1 _06111_ (
    .A(_00328_),
    .B(_00390_),
    .C(_00391_),
    .Y(_00151_)
  );
  NAND2X1 _06112_ (
    .A( dbg_0.mem_start ),
    .B(_00248_),
    .Y(_00392_)
  );
  NOR2X1 _06113_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00392_),
    .Y( dbg_0.dbg_i2c_0.mem_burst_rd )
  );
  OAI21X1 _06114_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00392_),
    .C(_00196_),
    .Y(_00393_)
  );
  NAND2X1 _06115_ (
    .A( dbg_0.mem_state_1_ ),
    .B( dbg_0.mem_ctl_2_ ),
    .Y(_00394_)
  );
  NOR2X1 _06116_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00394_),
    .Y(_00395_)
  );
  OR2X1 _06117_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00394_),
    .Y(_00396_)
  );
  OAI21X1 _06118_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00394_),
    .C(_00198_),
    .Y(_00397_)
  );
  MUX2X1 _06119_ (
    .A(_00397_),
    .B( dbg_0.dbg_i2c_0.dbg_rd ),
    .S(_00393_),
    .Y(_00398_)
  );
  INVX1 _06120_ (
    .A(_00398_),
    .Y(_00127_)
  );
  AOI21X1 _06121_ (
    .A(_00195_),
    .B( dbg_0.dbg_addr_1_ ),
    .C( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00399_)
  );
  NOR2X1 _06122_ (
    .A( dbg_0.dbg_addr_3_ ),
    .B(_00260_),
    .Y(_00400_)
  );
  NAND2X1 _06123_ (
    .A(_00261_),
    .B(_00400_),
    .Y(_00401_)
  );
  NOR2X1 _06124_ (
    .A(_00399_),
    .B(_00401_),
    .Y(_00402_)
  );
  NAND2X1 _06125_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00402_),
    .Y(_00403_)
  );
  NOR2X1 _06126_ (
    .A(_00194_),
    .B(_00403_),
    .Y(_00404_)
  );
  AND2X1 _06127_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00404_),
    .Y( dbg_0.istep )
  );
  NOR2X1 _06128_ (
    .A( dbg_0.inc_step_0_ ),
    .B( dbg_0.istep ),
    .Y(_00405_)
  );
  INVX1 _06129_ (
    .A(_00405_),
    .Y(_00128_)
  );
  NOR2X1 _06130_ (
    .A(_00214_),
    .B(_00253_),
    .Y(_05677_)
  );
  NOR2X1 _06131_ (
    .A(_00215_),
    .B(_00253_),
    .Y(_05684_)
  );
  NOR2X1 _06132_ (
    .A(_00216_),
    .B(_00253_),
    .Y(_05685_)
  );
  NOR2X1 _06133_ (
    .A(_00217_),
    .B(_00253_),
    .Y(_05686_)
  );
  NOR2X1 _06134_ (
    .A(_00218_),
    .B(_00253_),
    .Y(_05687_)
  );
  NOR2X1 _06135_ (
    .A(_00219_),
    .B(_00253_),
    .Y(_05688_)
  );
  NOR2X1 _06136_ (
    .A(_00220_),
    .B(_00253_),
    .Y(_05689_)
  );
  NOR2X1 _06137_ (
    .A(_00221_),
    .B(_00253_),
    .Y(_05690_)
  );
  OAI22X1 _06138_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00222_),
    .C(_00254_),
    .D(_00214_),
    .Y(_05691_)
  );
  OAI22X1 _06139_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00223_),
    .C(_00254_),
    .D(_00215_),
    .Y(_05692_)
  );
  OAI22X1 _06140_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00224_),
    .C(_00254_),
    .D(_00216_),
    .Y(_05678_)
  );
  OAI22X1 _06141_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00225_),
    .C(_00254_),
    .D(_00217_),
    .Y(_05679_)
  );
  OAI22X1 _06142_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00226_),
    .C(_00254_),
    .D(_00218_),
    .Y(_05680_)
  );
  OAI22X1 _06143_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00227_),
    .C(_00254_),
    .D(_00219_),
    .Y(_05681_)
  );
  OAI22X1 _06144_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00228_),
    .C(_00254_),
    .D(_00220_),
    .Y(_05682_)
  );
  OAI22X1 _06145_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00229_),
    .C(_00254_),
    .D(_00221_),
    .Y(_05683_)
  );
  NOR2X1 _06146_ (
    .A(_00326_),
    .B(_00401_),
    .Y(_00406_)
  );
  NAND3X1 _06147_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B( dbg_0.dbg_din_2_ ),
    .C(_00406_),
    .Y(_00407_)
  );
  AOI21X1 _06148_ (
    .A( dbg_0.cpu_stat_2_ ),
    .B(_00407_),
    .C(_05695_),
    .Y(_00408_)
  );
  INVX1 _06149_ (
    .A(_00408_),
    .Y(_00125_)
  );
  NAND3X1 _06150_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B( dbg_0.dbg_din_3_ ),
    .C(_00406_),
    .Y(_00409_)
  );
  NAND2X1 _06151_ (
    .A( dbg_0.cpu_stat_3_ ),
    .B(_00409_),
    .Y(_00410_)
  );
  NOR2X1 _06152_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B( dbg_0.fe_mdb_in_5_ ),
    .Y(_00411_)
  );
  NOR2X1 _06153_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .B( dbg_0.fe_mdb_in_4_ ),
    .Y(_00412_)
  );
  NAND3X1 _06154_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B( dbg_0.fe_mdb_in_0_ ),
    .C(_00412_),
    .Y(_00413_)
  );
  INVX1 _06155_ (
    .A(_00413_),
    .Y(_00414_)
  );
  NOR2X1 _06156_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_00202_),
    .Y(_00415_)
  );
  NAND3X1 _06157_ (
    .A( dbg_0.decode_noirq ),
    .B( dbg_0.cpu_ctl_3_ ),
    .C(_00415_),
    .Y(_00416_)
  );
  NOR2X1 _06158_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B( dbg_0.fe_mdb_in_12_ ),
    .Y(_00417_)
  );
  NOR2X1 _06159_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B( dbg_0.fe_mdb_in_10_ ),
    .Y(_00418_)
  );
  NAND2X1 _06160_ (
    .A(_00201_),
    .B( dbg_0.fe_mdb_in_6_ ),
    .Y(_00419_)
  );
  NAND2X1 _06161_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B( dbg_0.fe_mdb_in_8_ ),
    .Y(_00420_)
  );
  NOR2X1 _06162_ (
    .A(_00419_),
    .B(_00420_),
    .Y(_00421_)
  );
  NAND3X1 _06163_ (
    .A(_00417_),
    .B(_00418_),
    .C(_00421_),
    .Y(_00422_)
  );
  NOR2X1 _06164_ (
    .A(_00416_),
    .B(_00422_),
    .Y(_00423_)
  );
  NAND3X1 _06165_ (
    .A(_00411_),
    .B(_00414_),
    .C(_00423_),
    .Y(_00424_)
  );
  NAND2X1 _06166_ (
    .A(_00410_),
    .B(_00424_),
    .Y(_00126_)
  );
  NAND2X1 _06167_ (
    .A(_00195_),
    .B(_00258_),
    .Y(_00425_)
  );
  NOR2X1 _06168_ (
    .A(_00263_),
    .B(_00425_),
    .Y(_00426_)
  );
  NAND2X1 _06169_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00426_),
    .Y(_00427_)
  );
  NOR2X1 _06170_ (
    .A(_00200_),
    .B(_00427_),
    .Y(_00161_)
  );
  NOR2X1 _06171_ (
    .A(_00263_),
    .B(_00399_),
    .Y(_00428_)
  );
  NOR2X1 _06172_ (
    .A(_00259_),
    .B(_00401_),
    .Y(_00429_)
  );
  NOR2X1 _06173_ (
    .A(_00401_),
    .B(_00425_),
    .Y(_00430_)
  );
  NAND2X1 _06174_ (
    .A( dbg_0.dbg_addr_3_ ),
    .B( dbg_0.dbg_addr_4_ ),
    .Y(_00431_)
  );
  NOR2X1 _06175_ (
    .A( dbg_0.dbg_addr_5_ ),
    .B(_00431_),
    .Y(_00432_)
  );
  NAND2X1 _06176_ (
    .A(_00261_),
    .B(_00432_),
    .Y(_00433_)
  );
  NOR2X1 _06177_ (
    .A(_00425_),
    .B(_00433_),
    .Y(_00434_)
  );
  AOI22X1 _06178_ (
    .A( dbg_0.mem_cnt_0_ ),
    .B(_00327_),
    .C(_00429_),
    .D(1'h1),
    .Y(_00435_)
  );
  AOI22X1 _06179_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_00406_),
    .C(_00430_),
    .D(1'h1),
    .Y(_00436_)
  );
  INVX1 _06180_ (
    .A(_00436_),
    .Y(_00437_)
  );
  AOI21X1 _06181_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00437_),
    .Y(_00438_)
  );
  AOI22X1 _06182_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .B(_00264_),
    .C(_00428_),
    .D( dbg_0.mem_data_0_ ),
    .Y(_00439_)
  );
  NAND3X1 _06183_ (
    .A(_00435_),
    .B(_00438_),
    .C(_00439_),
    .Y( dbg_0.dbg_dout_0_ )
  );
  AOI22X1 _06184_ (
    .A( dbg_0.mem_data_1_ ),
    .B(_00428_),
    .C(_00429_),
    .D(1'h0),
    .Y(_00440_)
  );
  INVX1 _06185_ (
    .A(_00440_),
    .Y(_00441_)
  );
  AOI21X1 _06186_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .B(_00264_),
    .C(_00441_),
    .Y(_00442_)
  );
  AOI22X1 _06187_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00426_),
    .C(_00430_),
    .D(1'h1),
    .Y(_00443_)
  );
  AOI22X1 _06188_ (
    .A( dbg_0.mem_cnt_1_ ),
    .B(_00327_),
    .C(_00434_),
    .D(1'h0),
    .Y(_00444_)
  );
  NAND3X1 _06189_ (
    .A(_00442_),
    .B(_00443_),
    .C(_00444_),
    .Y( dbg_0.dbg_dout_1_ )
  );
  AOI22X1 _06190_ (
    .A( dbg_0.mem_cnt_2_ ),
    .B(_00327_),
    .C(_00428_),
    .D( dbg_0.mem_data_2_ ),
    .Y(_00445_)
  );
  INVX1 _06191_ (
    .A(_00445_),
    .Y(_00446_)
  );
  AOI21X1 _06192_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00446_),
    .Y(_00447_)
  );
  AOI22X1 _06193_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_00264_),
    .C(_00426_),
    .D( dbg_0.mem_ctl_2_ ),
    .Y(_00448_)
  );
  AOI22X1 _06194_ (
    .A( dbg_0.cpu_stat_2_ ),
    .B(_00406_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00449_)
  );
  INVX1 _06195_ (
    .A(_00449_),
    .Y(_00450_)
  );
  AOI21X1 _06196_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00450_),
    .Y(_00451_)
  );
  NAND3X1 _06197_ (
    .A(_00447_),
    .B(_00448_),
    .C(_00451_),
    .Y( dbg_0.dbg_dout_2_ )
  );
  AOI22X1 _06198_ (
    .A( dbg_0.cpu_ctl_3_ ),
    .B(_00402_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00452_)
  );
  AOI22X1 _06199_ (
    .A( dbg_0.mem_data_3_ ),
    .B(_00428_),
    .C(_00434_),
    .D(1'h0),
    .Y(_00453_)
  );
  AOI22X1 _06200_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_3_ ),
    .Y(_00454_)
  );
  NAND2X1 _06201_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00426_),
    .Y(_00455_)
  );
  AOI22X1 _06202_ (
    .A( dbg_0.cpu_stat_3_ ),
    .B(_00406_),
    .C(_00429_),
    .D(1'h0),
    .Y(_00456_)
  );
  NAND3X1 _06203_ (
    .A(_00454_),
    .B(_00455_),
    .C(_00456_),
    .Y(_00457_)
  );
  INVX1 _06204_ (
    .A(_00457_),
    .Y(_00458_)
  );
  NAND3X1 _06205_ (
    .A(_00452_),
    .B(_00453_),
    .C(_00458_),
    .Y( dbg_0.dbg_dout_3_ )
  );
  AOI22X1 _06206_ (
    .A( dbg_0.mem_data_4_ ),
    .B(_00428_),
    .C(_00434_),
    .D(1'h0),
    .Y(_00459_)
  );
  AOI22X1 _06207_ (
    .A( dbg_0.mem_cnt_4_ ),
    .B(_00327_),
    .C(_00402_),
    .D( dbg_0.cpu_ctl_4_ ),
    .Y(_00460_)
  );
  INVX1 _06208_ (
    .A(_00460_),
    .Y(_00461_)
  );
  AOI21X1 _06209_ (
    .A(1'h0),
    .B(_00430_),
    .C(_00461_),
    .Y(_00462_)
  );
  AOI22X1 _06210_ (
    .A( dbg_0.dbg_mem_addr_4_ ),
    .B(_00264_),
    .C(_00429_),
    .D(1'h0),
    .Y(_00463_)
  );
  NAND3X1 _06211_ (
    .A(_00459_),
    .B(_00462_),
    .C(_00463_),
    .Y( dbg_0.dbg_dout_4_ )
  );
  AOI22X1 _06212_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .B(_00264_),
    .C(_00402_),
    .D( dbg_0.cpu_ctl_5_ ),
    .Y(_00464_)
  );
  INVX1 _06213_ (
    .A(_00464_),
    .Y(_00465_)
  );
  AOI21X1 _06214_ (
    .A( dbg_0.mem_cnt_5_ ),
    .B(_00327_),
    .C(_00465_),
    .Y(_00466_)
  );
  AOI22X1 _06215_ (
    .A(1'h0),
    .B(_00430_),
    .C(_00434_),
    .D(1'h0),
    .Y(_00467_)
  );
  AOI22X1 _06216_ (
    .A( dbg_0.mem_data_5_ ),
    .B(_00428_),
    .C(_00429_),
    .D(1'h0),
    .Y(_00468_)
  );
  NAND3X1 _06217_ (
    .A(_00466_),
    .B(_00467_),
    .C(_00468_),
    .Y( dbg_0.dbg_dout_5_ )
  );
  AOI22X1 _06218_ (
    .A( clock_module_0.dbg_cpu_reset ),
    .B(_00402_),
    .C(_00429_),
    .D(1'h0),
    .Y(_00469_)
  );
  INVX1 _06219_ (
    .A(_00469_),
    .Y(_00470_)
  );
  AOI22X1 _06220_ (
    .A( dbg_0.mem_cnt_6_ ),
    .B(_00327_),
    .C(_00428_),
    .D( dbg_0.mem_data_6_ ),
    .Y(_00471_)
  );
  AOI21X1 _06221_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00470_),
    .Y(_00472_)
  );
  AOI22X1 _06222_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .B(_00264_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00473_)
  );
  NAND3X1 _06223_ (
    .A(_00471_),
    .B(_00472_),
    .C(_00473_),
    .Y( dbg_0.dbg_dout_6_ )
  );
  AOI22X1 _06224_ (
    .A( dbg_0.dbg_mem_addr_7_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_7_ ),
    .Y(_00474_)
  );
  NAND2X1 _06225_ (
    .A( dbg_0.mem_data_7_ ),
    .B(_00428_),
    .Y(_00475_)
  );
  AOI22X1 _06226_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00476_)
  );
  INVX1 _06227_ (
    .A(_00476_),
    .Y(_00477_)
  );
  AOI21X1 _06228_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00477_),
    .Y(_00478_)
  );
  NAND3X1 _06229_ (
    .A(_00474_),
    .B(_00475_),
    .C(_00478_),
    .Y( dbg_0.dbg_dout_7_ )
  );
  AOI22X1 _06230_ (
    .A( dbg_0.dbg_mem_addr_8_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_8_ ),
    .Y(_00479_)
  );
  NAND2X1 _06231_ (
    .A( dbg_0.mem_data_8_ ),
    .B(_00428_),
    .Y(_00480_)
  );
  AOI22X1 _06232_ (
    .A(1'h1),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00481_)
  );
  INVX1 _06233_ (
    .A(_00481_),
    .Y(_00482_)
  );
  AOI21X1 _06234_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00482_),
    .Y(_00483_)
  );
  NAND3X1 _06235_ (
    .A(_00479_),
    .B(_00480_),
    .C(_00483_),
    .Y( dbg_0.dbg_dout_8_ )
  );
  AOI22X1 _06236_ (
    .A( dbg_0.dbg_mem_addr_9_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_9_ ),
    .Y(_00484_)
  );
  NAND2X1 _06237_ (
    .A(1'h0),
    .B(_00434_),
    .Y(_00485_)
  );
  AOI22X1 _06238_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00486_)
  );
  INVX1 _06239_ (
    .A(_00486_),
    .Y(_00487_)
  );
  AOI21X1 _06240_ (
    .A( dbg_0.mem_data_9_ ),
    .B(_00428_),
    .C(_00487_),
    .Y(_00488_)
  );
  NAND3X1 _06241_ (
    .A(_00484_),
    .B(_00485_),
    .C(_00488_),
    .Y( dbg_0.dbg_dout_9_ )
  );
  AOI22X1 _06242_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_10_ ),
    .Y(_00489_)
  );
  NAND2X1 _06243_ (
    .A(1'h0),
    .B(_00434_),
    .Y(_00490_)
  );
  AOI22X1 _06244_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00491_)
  );
  INVX1 _06245_ (
    .A(_00491_),
    .Y(_00492_)
  );
  AOI21X1 _06246_ (
    .A( dbg_0.mem_data_10_ ),
    .B(_00428_),
    .C(_00492_),
    .Y(_00493_)
  );
  NAND3X1 _06247_ (
    .A(_00489_),
    .B(_00490_),
    .C(_00493_),
    .Y( dbg_0.dbg_dout_10_ )
  );
  AOI22X1 _06248_ (
    .A( dbg_0.dbg_mem_addr_11_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_11_ ),
    .Y(_00494_)
  );
  NAND2X1 _06249_ (
    .A( dbg_0.mem_data_11_ ),
    .B(_00428_),
    .Y(_00495_)
  );
  AOI22X1 _06250_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00496_)
  );
  INVX1 _06251_ (
    .A(_00496_),
    .Y(_00497_)
  );
  AOI21X1 _06252_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00497_),
    .Y(_00498_)
  );
  NAND3X1 _06253_ (
    .A(_00494_),
    .B(_00495_),
    .C(_00498_),
    .Y( dbg_0.dbg_dout_11_ )
  );
  NAND2X1 _06254_ (
    .A( dbg_0.mem_data_12_ ),
    .B(_00428_),
    .Y(_00499_)
  );
  AOI22X1 _06255_ (
    .A( dbg_0.dbg_mem_addr_12_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_12_ ),
    .Y(_00500_)
  );
  INVX1 _06256_ (
    .A(_00500_),
    .Y(_00501_)
  );
  AOI22X1 _06257_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00502_)
  );
  AOI21X1 _06258_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00501_),
    .Y(_00503_)
  );
  NAND3X1 _06259_ (
    .A(_00499_),
    .B(_00502_),
    .C(_00503_),
    .Y( dbg_0.dbg_dout_12_ )
  );
  AOI22X1 _06260_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_13_ ),
    .Y(_00504_)
  );
  NAND2X1 _06261_ (
    .A(1'h0),
    .B(_00434_),
    .Y(_00505_)
  );
  AOI22X1 _06262_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h0),
    .Y(_00506_)
  );
  INVX1 _06263_ (
    .A(_00506_),
    .Y(_00507_)
  );
  AOI21X1 _06264_ (
    .A( dbg_0.mem_data_13_ ),
    .B(_00428_),
    .C(_00507_),
    .Y(_00508_)
  );
  NAND3X1 _06265_ (
    .A(_00504_),
    .B(_00505_),
    .C(_00508_),
    .Y( dbg_0.dbg_dout_13_ )
  );
  NAND2X1 _06266_ (
    .A( dbg_0.mem_data_14_ ),
    .B(_00428_),
    .Y(_00509_)
  );
  AOI22X1 _06267_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_14_ ),
    .Y(_00510_)
  );
  INVX1 _06268_ (
    .A(_00510_),
    .Y(_00511_)
  );
  AOI22X1 _06269_ (
    .A(1'h0),
    .B(_00429_),
    .C(_00430_),
    .D(1'h1),
    .Y(_00512_)
  );
  AOI21X1 _06270_ (
    .A(1'h0),
    .B(_00434_),
    .C(_00511_),
    .Y(_00513_)
  );
  NAND3X1 _06271_ (
    .A(_00509_),
    .B(_00512_),
    .C(_00513_),
    .Y( dbg_0.dbg_dout_14_ )
  );
  AOI22X1 _06272_ (
    .A(1'h1),
    .B(_00429_),
    .C(_00434_),
    .D(1'h0),
    .Y(_00514_)
  );
  INVX1 _06273_ (
    .A(_00514_),
    .Y(_00515_)
  );
  AOI21X1 _06274_ (
    .A( dbg_0.mem_data_15_ ),
    .B(_00428_),
    .C(_00515_),
    .Y(_00516_)
  );
  NAND2X1 _06275_ (
    .A(1'h0),
    .B(_00430_),
    .Y(_00517_)
  );
  AOI22X1 _06276_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .B(_00264_),
    .C(_00327_),
    .D( dbg_0.mem_cnt_15_ ),
    .Y(_00518_)
  );
  NAND3X1 _06277_ (
    .A(_00516_),
    .B(_00517_),
    .C(_00518_),
    .Y( dbg_0.dbg_dout_15_ )
  );
  OAI21X1 _06278_ (
    .A( dbg_0.cpu_ctl_4_ ),
    .B(_00230_),
    .C( dbg_0.cpu_stat_full_0_ ),
    .Y(_00519_)
  );
  INVX1 _06279_ (
    .A(_00519_),
    .Y(_05582_)
  );
  OAI22X1 _06280_ (
    .A( dbg_0.mem_state_0_ ),
    .B(_00251_),
    .C(_00403_),
    .D(_00200_),
    .Y(_00520_)
  );
  AND2X1 _06281_ (
    .A( dbg_0.cpu_ctl_5_ ),
    .B(_05695_),
    .Y(_00521_)
  );
  AOI21X1 _06282_ (
    .A(dbg_en),
    .B(_00521_),
    .C( dbg_0.halt_flag ),
    .Y(_00522_)
  );
  NAND2X1 _06283_ (
    .A(_00424_),
    .B(_00522_),
    .Y(_00523_)
  );
  AOI21X1 _06284_ (
    .A(_00194_),
    .B(_00520_),
    .C(_00523_),
    .Y(_00524_)
  );
  NOR2X1 _06285_ (
    .A( dbg_0.inc_step_1_ ),
    .B(_00524_),
    .Y( dbg_0.dbg_halt_cmd )
  );
  NOR2X1 _06286_ (
    .A(_00197_),
    .B(_00392_),
    .Y( dbg_0.dbg_i2c_0.mem_burst_wr )
  );
  OAI21X1 _06287_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B( dbg_0.dbg_i2c_0.dbg_rd ),
    .C( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00525_)
  );
  OAI21X1 _06288_ (
    .A( dbg_0.mem_ctl_1_ ),
    .B(_00392_),
    .C(_00525_),
    .Y(_00162_)
  );
  AND2X1 _06289_ (
    .A(_00197_),
    .B( dbg_0.dbg_mem_en ),
    .Y( dbg_0.dbg_mem_rd )
  );
  MUX2X1 _06290_ (
    .A( dbg_0.cpu_ctl_3_ ),
    .B( dbg_0.dbg_din_3_ ),
    .S(_00403_),
    .Y(_00526_)
  );
  INVX1 _06291_ (
    .A(_00526_),
    .Y(_00164_)
  );
  MUX2X1 _06292_ (
    .A( dbg_0.cpu_ctl_4_ ),
    .B( dbg_0.dbg_din_4_ ),
    .S(_00403_),
    .Y(_00527_)
  );
  INVX1 _06293_ (
    .A(_00527_),
    .Y(_00165_)
  );
  MUX2X1 _06294_ (
    .A( dbg_0.cpu_ctl_5_ ),
    .B( dbg_0.dbg_din_5_ ),
    .S(_00403_),
    .Y(_00528_)
  );
  INVX1 _06295_ (
    .A(_00528_),
    .Y(_00166_)
  );
  MUX2X1 _06296_ (
    .A( clock_module_0.dbg_cpu_reset ),
    .B( dbg_0.dbg_din_6_ ),
    .S(_00403_),
    .Y(_00529_)
  );
  INVX1 _06297_ (
    .A(_00529_),
    .Y(_00167_)
  );
  AOI21X1 _06298_ (
    .A(_00196_),
    .B(_00392_),
    .C( dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00168_)
  );
  NAND2X1 _06299_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00404_),
    .Y(_00530_)
  );
  OAI21X1 _06300_ (
    .A(_00193_),
    .B( dbg_0.mem_state_0_ ),
    .C(_00530_),
    .Y(_00531_)
  );
  NOR2X1 _06301_ (
    .A(_00524_),
    .B(_00531_),
    .Y(_00169_)
  );
  NAND2X1 _06302_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00428_),
    .Y(_00532_)
  );
  AOI21X1 _06303_ (
    .A( dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00428_),
    .C(_00397_),
    .Y(_00533_)
  );
  NAND3X1 _06304_ (
    .A(_00198_),
    .B(_00396_),
    .C(_00532_),
    .Y(_00534_)
  );
  MUX2X1 _06305_ (
    .A( dbg_0.dbg_mem_din_0_ ),
    .B( dbg_0.dbg_mem_din_8_ ),
    .S(_00254_),
    .Y(_00535_)
  );
  AND2X1 _06306_ (
    .A(_00396_),
    .B(_00535_),
    .Y(_00536_)
  );
  OAI21X1 _06307_ (
    .A( dbg_0.dbg_reg_din_0_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00537_)
  );
  OAI21X1 _06308_ (
    .A(_00536_),
    .B(_00537_),
    .C(_00532_),
    .Y(_00538_)
  );
  OAI21X1 _06309_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00532_),
    .C(_00538_),
    .Y(_00539_)
  );
  OAI21X1 _06310_ (
    .A(_00214_),
    .B(_00534_),
    .C(_00539_),
    .Y(_00170_)
  );
  MUX2X1 _06311_ (
    .A( dbg_0.dbg_mem_din_1_ ),
    .B( dbg_0.dbg_mem_din_9_ ),
    .S(_00254_),
    .Y(_00540_)
  );
  AND2X1 _06312_ (
    .A(_00396_),
    .B(_00540_),
    .Y(_00541_)
  );
  OAI21X1 _06313_ (
    .A( dbg_0.dbg_reg_din_1_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00542_)
  );
  OAI21X1 _06314_ (
    .A(_00541_),
    .B(_00542_),
    .C(_00532_),
    .Y(_00543_)
  );
  OAI21X1 _06315_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00532_),
    .C(_00543_),
    .Y(_00544_)
  );
  OAI21X1 _06316_ (
    .A(_00215_),
    .B(_00534_),
    .C(_00544_),
    .Y(_00171_)
  );
  MUX2X1 _06317_ (
    .A( dbg_0.dbg_mem_din_2_ ),
    .B( dbg_0.dbg_mem_din_10_ ),
    .S(_00254_),
    .Y(_00545_)
  );
  AND2X1 _06318_ (
    .A(_00396_),
    .B(_00545_),
    .Y(_00546_)
  );
  OAI21X1 _06319_ (
    .A( dbg_0.dbg_reg_din_2_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00547_)
  );
  OAI21X1 _06320_ (
    .A(_00546_),
    .B(_00547_),
    .C(_00532_),
    .Y(_00548_)
  );
  OAI21X1 _06321_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00532_),
    .C(_00548_),
    .Y(_00549_)
  );
  OAI21X1 _06322_ (
    .A(_00216_),
    .B(_00534_),
    .C(_00549_),
    .Y(_00172_)
  );
  MUX2X1 _06323_ (
    .A( dbg_0.dbg_mem_din_3_ ),
    .B( dbg_0.dbg_mem_din_11_ ),
    .S(_00254_),
    .Y(_00550_)
  );
  AND2X1 _06324_ (
    .A(_00396_),
    .B(_00550_),
    .Y(_00551_)
  );
  OAI21X1 _06325_ (
    .A( dbg_0.dbg_reg_din_3_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00552_)
  );
  OAI21X1 _06326_ (
    .A(_00551_),
    .B(_00552_),
    .C(_00532_),
    .Y(_00553_)
  );
  OAI21X1 _06327_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00532_),
    .C(_00553_),
    .Y(_00554_)
  );
  OAI21X1 _06328_ (
    .A(_00217_),
    .B(_00534_),
    .C(_00554_),
    .Y(_00173_)
  );
  MUX2X1 _06329_ (
    .A( dbg_0.dbg_mem_din_4_ ),
    .B( dbg_0.dbg_mem_din_12_ ),
    .S(_00254_),
    .Y(_00555_)
  );
  AND2X1 _06330_ (
    .A(_00396_),
    .B(_00555_),
    .Y(_00556_)
  );
  OAI21X1 _06331_ (
    .A( dbg_0.dbg_reg_din_4_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00557_)
  );
  OAI21X1 _06332_ (
    .A(_00556_),
    .B(_00557_),
    .C(_00532_),
    .Y(_00558_)
  );
  OAI21X1 _06333_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00532_),
    .C(_00558_),
    .Y(_00559_)
  );
  OAI21X1 _06334_ (
    .A(_00218_),
    .B(_00534_),
    .C(_00559_),
    .Y(_00174_)
  );
  MUX2X1 _06335_ (
    .A( dbg_0.dbg_mem_din_5_ ),
    .B( dbg_0.dbg_mem_din_13_ ),
    .S(_00254_),
    .Y(_00560_)
  );
  AND2X1 _06336_ (
    .A(_00396_),
    .B(_00560_),
    .Y(_00561_)
  );
  OAI21X1 _06337_ (
    .A( dbg_0.dbg_reg_din_5_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00562_)
  );
  OAI21X1 _06338_ (
    .A(_00561_),
    .B(_00562_),
    .C(_00532_),
    .Y(_00563_)
  );
  OAI21X1 _06339_ (
    .A( dbg_0.dbg_din_5_ ),
    .B(_00532_),
    .C(_00563_),
    .Y(_00564_)
  );
  OAI21X1 _06340_ (
    .A(_00219_),
    .B(_00534_),
    .C(_00564_),
    .Y(_00175_)
  );
  MUX2X1 _06341_ (
    .A( dbg_0.dbg_mem_din_6_ ),
    .B( dbg_0.dbg_mem_din_14_ ),
    .S(_00254_),
    .Y(_00565_)
  );
  AND2X1 _06342_ (
    .A(_00396_),
    .B(_00565_),
    .Y(_00566_)
  );
  OAI21X1 _06343_ (
    .A( dbg_0.dbg_reg_din_6_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00567_)
  );
  OAI21X1 _06344_ (
    .A(_00566_),
    .B(_00567_),
    .C(_00532_),
    .Y(_00568_)
  );
  OAI21X1 _06345_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00532_),
    .C(_00568_),
    .Y(_00569_)
  );
  OAI21X1 _06346_ (
    .A(_00220_),
    .B(_00534_),
    .C(_00569_),
    .Y(_00176_)
  );
  MUX2X1 _06347_ (
    .A( dbg_0.dbg_mem_din_7_ ),
    .B( dbg_0.dbg_mem_din_15_ ),
    .S(_00254_),
    .Y(_00570_)
  );
  AND2X1 _06348_ (
    .A(_00396_),
    .B(_00570_),
    .Y(_00571_)
  );
  OAI21X1 _06349_ (
    .A( dbg_0.dbg_reg_din_7_ ),
    .B(_00396_),
    .C(_00397_),
    .Y(_00572_)
  );
  OAI21X1 _06350_ (
    .A(_00571_),
    .B(_00572_),
    .C(_00532_),
    .Y(_00573_)
  );
  OAI21X1 _06351_ (
    .A( dbg_0.dbg_din_7_ ),
    .B(_00532_),
    .C(_00573_),
    .Y(_00574_)
  );
  OAI21X1 _06352_ (
    .A(_00221_),
    .B(_00534_),
    .C(_00574_),
    .Y(_00177_)
  );
  NAND2X1 _06353_ (
    .A( dbg_0.dbg_reg_din_8_ ),
    .B(_00395_),
    .Y(_00575_)
  );
  NOR2X1 _06354_ (
    .A(_00198_),
    .B( dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00576_)
  );
  NAND2X1 _06355_ (
    .A( dbg_0.dbg_mem_din_8_ ),
    .B(_00576_),
    .Y(_00577_)
  );
  OAI21X1 _06356_ (
    .A(_00395_),
    .B(_00577_),
    .C(_00575_),
    .Y(_00578_)
  );
  AOI22X1 _06357_ (
    .A( dbg_0.mem_data_8_ ),
    .B(_00533_),
    .C(_00578_),
    .D(_00532_),
    .Y(_00579_)
  );
  OAI21X1 _06358_ (
    .A(_00208_),
    .B(_00532_),
    .C(_00579_),
    .Y(_00178_)
  );
  NAND2X1 _06359_ (
    .A( dbg_0.dbg_reg_din_9_ ),
    .B(_00395_),
    .Y(_00580_)
  );
  NAND2X1 _06360_ (
    .A( dbg_0.dbg_mem_din_9_ ),
    .B(_00576_),
    .Y(_00581_)
  );
  OAI21X1 _06361_ (
    .A(_00395_),
    .B(_00581_),
    .C(_00580_),
    .Y(_00582_)
  );
  AOI22X1 _06362_ (
    .A( dbg_0.mem_data_9_ ),
    .B(_00533_),
    .C(_00582_),
    .D(_00532_),
    .Y(_00583_)
  );
  OAI21X1 _06363_ (
    .A(_00210_),
    .B(_00532_),
    .C(_00583_),
    .Y(_00179_)
  );
  NAND2X1 _06364_ (
    .A( dbg_0.dbg_reg_din_10_ ),
    .B(_00395_),
    .Y(_00584_)
  );
  NAND2X1 _06365_ (
    .A( dbg_0.dbg_mem_din_10_ ),
    .B(_00576_),
    .Y(_00585_)
  );
  OAI21X1 _06366_ (
    .A(_00395_),
    .B(_00585_),
    .C(_00584_),
    .Y(_00586_)
  );
  MUX2X1 _06367_ (
    .A(_00586_),
    .B( dbg_0.dbg_din_10_ ),
    .S(_00532_),
    .Y(_00587_)
  );
  OAI21X1 _06368_ (
    .A(_00224_),
    .B(_00534_),
    .C(_00587_),
    .Y(_00180_)
  );
  NAND2X1 _06369_ (
    .A( dbg_0.dbg_reg_din_11_ ),
    .B(_00395_),
    .Y(_00588_)
  );
  NAND2X1 _06370_ (
    .A( dbg_0.dbg_mem_din_11_ ),
    .B(_00576_),
    .Y(_00589_)
  );
  OAI21X1 _06371_ (
    .A(_00395_),
    .B(_00589_),
    .C(_00588_),
    .Y(_00590_)
  );
  MUX2X1 _06372_ (
    .A(_00590_),
    .B( dbg_0.dbg_din_11_ ),
    .S(_00532_),
    .Y(_00591_)
  );
  OAI21X1 _06373_ (
    .A(_00225_),
    .B(_00534_),
    .C(_00591_),
    .Y(_00181_)
  );
  NAND2X1 _06374_ (
    .A( dbg_0.dbg_reg_din_12_ ),
    .B(_00395_),
    .Y(_00592_)
  );
  NAND2X1 _06375_ (
    .A( dbg_0.dbg_mem_din_12_ ),
    .B(_00576_),
    .Y(_00593_)
  );
  OAI21X1 _06376_ (
    .A(_00395_),
    .B(_00593_),
    .C(_00592_),
    .Y(_00594_)
  );
  MUX2X1 _06377_ (
    .A(_00594_),
    .B( dbg_0.dbg_din_12_ ),
    .S(_00532_),
    .Y(_00595_)
  );
  OAI21X1 _06378_ (
    .A(_00226_),
    .B(_00534_),
    .C(_00595_),
    .Y(_00182_)
  );
  NAND2X1 _06379_ (
    .A( dbg_0.dbg_reg_din_13_ ),
    .B(_00395_),
    .Y(_00596_)
  );
  NAND2X1 _06380_ (
    .A( dbg_0.dbg_mem_din_13_ ),
    .B(_00576_),
    .Y(_00597_)
  );
  OAI21X1 _06381_ (
    .A(_00395_),
    .B(_00597_),
    .C(_00596_),
    .Y(_00598_)
  );
  AOI22X1 _06382_ (
    .A( dbg_0.mem_data_13_ ),
    .B(_00533_),
    .C(_00598_),
    .D(_00532_),
    .Y(_00599_)
  );
  OAI21X1 _06383_ (
    .A(_00212_),
    .B(_00532_),
    .C(_00599_),
    .Y(_00183_)
  );
  NAND2X1 _06384_ (
    .A( dbg_0.dbg_reg_din_14_ ),
    .B(_00395_),
    .Y(_00600_)
  );
  NAND2X1 _06385_ (
    .A( dbg_0.dbg_mem_din_14_ ),
    .B(_00576_),
    .Y(_00601_)
  );
  OAI21X1 _06386_ (
    .A(_00395_),
    .B(_00601_),
    .C(_00600_),
    .Y(_00602_)
  );
  MUX2X1 _06387_ (
    .A(_00602_),
    .B( dbg_0.dbg_din_14_ ),
    .S(_00532_),
    .Y(_00603_)
  );
  OAI21X1 _06388_ (
    .A(_00228_),
    .B(_00534_),
    .C(_00603_),
    .Y(_00184_)
  );
  NAND2X1 _06389_ (
    .A( dbg_0.dbg_reg_din_15_ ),
    .B(_00395_),
    .Y(_00604_)
  );
  NAND2X1 _06390_ (
    .A( dbg_0.dbg_mem_din_15_ ),
    .B(_00576_),
    .Y(_00605_)
  );
  OAI21X1 _06391_ (
    .A(_00395_),
    .B(_00605_),
    .C(_00604_),
    .Y(_00606_)
  );
  AOI22X1 _06392_ (
    .A( dbg_0.mem_data_15_ ),
    .B(_00533_),
    .C(_00606_),
    .D(_00532_),
    .Y(_00607_)
  );
  OAI21X1 _06393_ (
    .A(_00213_),
    .B(_00532_),
    .C(_00607_),
    .Y(_00185_)
  );
  NAND2X1 _06394_ (
    .A(_00197_),
    .B(_00427_),
    .Y(_00608_)
  );
  OAI21X1 _06395_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00427_),
    .C(_00608_),
    .Y(_00609_)
  );
  INVX1 _06396_ (
    .A(_00609_),
    .Y(_00186_)
  );
  MUX2X1 _06397_ (
    .A( dbg_0.mem_ctl_2_ ),
    .B( dbg_0.dbg_din_2_ ),
    .S(_00427_),
    .Y(_00610_)
  );
  INVX1 _06398_ (
    .A(_00610_),
    .Y(_00187_)
  );
  MUX2X1 _06399_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .B( dbg_0.dbg_din_3_ ),
    .S(_00427_),
    .Y(_00611_)
  );
  INVX1 _06400_ (
    .A(_00611_),
    .Y(_00188_)
  );
  DFFSR _06401_ (
    .CLK(dco_clk),
    .D(_00164_),
    .Q( dbg_0.cpu_ctl_3_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06402_ (
    .CLK(dco_clk),
    .D(_00165_),
    .Q( dbg_0.cpu_ctl_4_ ),
    .R(1'h1),
    .S(_00163_)
  );
  DFFSR _06403_ (
    .CLK(dco_clk),
    .D(_00166_),
    .Q( dbg_0.cpu_ctl_5_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06404_ (
    .CLK(dco_clk),
    .D(_00167_),
    .Q( clock_module_0.dbg_cpu_reset ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06405_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_mem_rd ),
    .Q( dbg_0.dbg_mem_rd_dly ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06406_ (
    .CLK(dco_clk),
    .D( dbg_0.mem_state_nxt_0_ ),
    .Q( dbg_0.mem_state_0_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06407_ (
    .CLK(dco_clk),
    .D( dbg_0.mem_state_nxt_1_ ),
    .Q( dbg_0.mem_state_1_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06408_ (
    .CLK(dco_clk),
    .D(_00162_),
    .Q( dbg_0.mem_startb ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06409_ (
    .CLK(dco_clk),
    .D(_00168_),
    .Q( dbg_0.dbg_i2c_0.mem_burst ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06410_ (
    .CLK(dco_clk),
    .D( dbg_0.istep ),
    .Q( dbg_0.inc_step_0_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06411_ (
    .CLK(dco_clk),
    .D(_00128_),
    .Q( dbg_0.inc_step_1_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06412_ (
    .CLK(dco_clk),
    .D(_00127_),
    .Q( dbg_0.dbg_rd_rdy ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06413_ (
    .CLK(dco_clk),
    .D(_00145_),
    .Q( dbg_0.mem_cnt_0_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06414_ (
    .CLK(dco_clk),
    .D(_00152_),
    .Q( dbg_0.mem_cnt_1_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06415_ (
    .CLK(dco_clk),
    .D(_00153_),
    .Q( dbg_0.mem_cnt_2_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06416_ (
    .CLK(dco_clk),
    .D(_00154_),
    .Q( dbg_0.mem_cnt_3_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06417_ (
    .CLK(dco_clk),
    .D(_00155_),
    .Q( dbg_0.mem_cnt_4_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06418_ (
    .CLK(dco_clk),
    .D(_00156_),
    .Q( dbg_0.mem_cnt_5_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06419_ (
    .CLK(dco_clk),
    .D(_00157_),
    .Q( dbg_0.mem_cnt_6_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06420_ (
    .CLK(dco_clk),
    .D(_00158_),
    .Q( dbg_0.mem_cnt_7_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06421_ (
    .CLK(dco_clk),
    .D(_00159_),
    .Q( dbg_0.mem_cnt_8_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06422_ (
    .CLK(dco_clk),
    .D(_00160_),
    .Q( dbg_0.mem_cnt_9_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06423_ (
    .CLK(dco_clk),
    .D(_00146_),
    .Q( dbg_0.mem_cnt_10_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06424_ (
    .CLK(dco_clk),
    .D(_00147_),
    .Q( dbg_0.mem_cnt_11_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06425_ (
    .CLK(dco_clk),
    .D(_00148_),
    .Q( dbg_0.mem_cnt_12_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06426_ (
    .CLK(dco_clk),
    .D(_00149_),
    .Q( dbg_0.mem_cnt_13_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06427_ (
    .CLK(dco_clk),
    .D(_00150_),
    .Q( dbg_0.mem_cnt_14_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06428_ (
    .CLK(dco_clk),
    .D(_00151_),
    .Q( dbg_0.mem_cnt_15_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06429_ (
    .CLK(dco_clk),
    .D(_00129_),
    .Q( dbg_0.dbg_mem_addr_0_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06430_ (
    .CLK(dco_clk),
    .D(_00136_),
    .Q( dbg_0.dbg_mem_addr_1_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06431_ (
    .CLK(dco_clk),
    .D(_00137_),
    .Q( dbg_0.dbg_mem_addr_2_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06432_ (
    .CLK(dco_clk),
    .D(_00138_),
    .Q( dbg_0.dbg_mem_addr_3_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06433_ (
    .CLK(dco_clk),
    .D(_00139_),
    .Q( dbg_0.dbg_mem_addr_4_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06434_ (
    .CLK(dco_clk),
    .D(_00140_),
    .Q( dbg_0.dbg_mem_addr_5_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06435_ (
    .CLK(dco_clk),
    .D(_00141_),
    .Q( dbg_0.dbg_mem_addr_6_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06436_ (
    .CLK(dco_clk),
    .D(_00142_),
    .Q( dbg_0.dbg_mem_addr_7_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06437_ (
    .CLK(dco_clk),
    .D(_00143_),
    .Q( dbg_0.dbg_mem_addr_8_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06438_ (
    .CLK(dco_clk),
    .D(_00144_),
    .Q( dbg_0.dbg_mem_addr_9_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06439_ (
    .CLK(dco_clk),
    .D(_00130_),
    .Q( dbg_0.dbg_mem_addr_10_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06440_ (
    .CLK(dco_clk),
    .D(_00131_),
    .Q( dbg_0.dbg_mem_addr_11_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06441_ (
    .CLK(dco_clk),
    .D(_00132_),
    .Q( dbg_0.dbg_mem_addr_12_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06442_ (
    .CLK(dco_clk),
    .D(_00133_),
    .Q( dbg_0.dbg_mem_addr_13_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06443_ (
    .CLK(dco_clk),
    .D(_00134_),
    .Q( dbg_0.dbg_mem_addr_14_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06444_ (
    .CLK(dco_clk),
    .D(_00135_),
    .Q( dbg_0.dbg_mem_addr_15_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06445_ (
    .CLK(dco_clk),
    .D(_00169_),
    .Q( dbg_0.halt_flag ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06446_ (
    .CLK(dco_clk),
    .D(_00161_),
    .Q( dbg_0.mem_start ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06447_ (
    .CLK(dco_clk),
    .D(_00170_),
    .Q( dbg_0.mem_data_0_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06448_ (
    .CLK(dco_clk),
    .D(_00171_),
    .Q( dbg_0.mem_data_1_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06449_ (
    .CLK(dco_clk),
    .D(_00172_),
    .Q( dbg_0.mem_data_2_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06450_ (
    .CLK(dco_clk),
    .D(_00173_),
    .Q( dbg_0.mem_data_3_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06451_ (
    .CLK(dco_clk),
    .D(_00174_),
    .Q( dbg_0.mem_data_4_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06452_ (
    .CLK(dco_clk),
    .D(_00175_),
    .Q( dbg_0.mem_data_5_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06453_ (
    .CLK(dco_clk),
    .D(_00176_),
    .Q( dbg_0.mem_data_6_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06454_ (
    .CLK(dco_clk),
    .D(_00177_),
    .Q( dbg_0.mem_data_7_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06455_ (
    .CLK(dco_clk),
    .D(_00178_),
    .Q( dbg_0.mem_data_8_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06456_ (
    .CLK(dco_clk),
    .D(_00179_),
    .Q( dbg_0.mem_data_9_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06457_ (
    .CLK(dco_clk),
    .D(_00180_),
    .Q( dbg_0.mem_data_10_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06458_ (
    .CLK(dco_clk),
    .D(_00181_),
    .Q( dbg_0.mem_data_11_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06459_ (
    .CLK(dco_clk),
    .D(_00182_),
    .Q( dbg_0.mem_data_12_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06460_ (
    .CLK(dco_clk),
    .D(_00183_),
    .Q( dbg_0.mem_data_13_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06461_ (
    .CLK(dco_clk),
    .D(_00184_),
    .Q( dbg_0.mem_data_14_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06462_ (
    .CLK(dco_clk),
    .D(_00185_),
    .Q( dbg_0.mem_data_15_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06463_ (
    .CLK(dco_clk),
    .D(_00125_),
    .Q( dbg_0.cpu_stat_2_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06464_ (
    .CLK(dco_clk),
    .D(_00126_),
    .Q( dbg_0.cpu_stat_3_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06465_ (
    .CLK(dco_clk),
    .D(_00186_),
    .Q( dbg_0.mem_ctl_1_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06466_ (
    .CLK(dco_clk),
    .D(_00187_),
    .Q( dbg_0.mem_ctl_2_ ),
    .R(_00163_),
    .S(1'h1)
  );
  DFFSR _06467_ (
    .CLK(dco_clk),
    .D(_00188_),
    .Q( dbg_0.dbg_i2c_0.mem_bw ),
    .R(_00163_),
    .S(1'h1)
  );
  INVX1 _06468_ (
    .A( dbg_0.dbg_i2c_0.scl_sync_n ),
    .Y( dbg_0.dbg_i2c_0.scl_sync )
  );
  INVX1 _06469_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .Y(_00649_)
  );
  INVX1 _06470_ (
    .A( dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .Y( dbg_0.dbg_i2c_0.sda_in_sync )
  );
  INVX1 _06471_ (
    .A( dbg_0.dbg_i2c_0.sda_in_dly ),
    .Y(_00650_)
  );
  INVX1 _06472_ (
    .A( dbg_0.dbg_i2c_0.i2c_active_seq ),
    .Y(_00651_)
  );
  INVX1 _06473_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .Y(_00652_)
  );
  INVX1 _06474_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00653_)
  );
  INVX1 _06475_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00654_)
  );
  INVX1 _06476_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .Y(_00655_)
  );
  INVX1 _06477_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .Y(_00656_)
  );
  INVX1 _06478_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .Y(_00657_)
  );
  INVX1 _06479_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .Y(_00658_)
  );
  INVX1 _06480_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .Y(_00659_)
  );
  INVX1 _06481_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00660_)
  );
  INVX1 _06482_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .Y(_00661_)
  );
  INVX1 _06483_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00662_)
  );
  INVX1 _06484_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .Y(_00663_)
  );
  INVX1 _06485_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .Y(_00664_)
  );
  INVX1 _06486_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00665_)
  );
  INVX1 _06487_ (
    .A( dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00666_)
  );
  INVX1 _06488_ (
    .A(dbg_i2c_scl),
    .Y( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in )
  );
  INVX1 _06489_ (
    .A(dbg_i2c_sda_in),
    .Y( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in )
  );
  INVX1 _06490_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00614_)
  );
  INVX1 _06491_ (
    .A( dbg_0.dbg_din_11_ ),
    .Y(_00667_)
  );
  INVX1 _06492_ (
    .A( dbg_0.dbg_din_12_ ),
    .Y(_00668_)
  );
  INVX1 _06493_ (
    .A( dbg_0.dbg_din_13_ ),
    .Y(_00669_)
  );
  INVX1 _06494_ (
    .A( dbg_0.dbg_din_14_ ),
    .Y(_00670_)
  );
  INVX1 _06495_ (
    .A( dbg_0.dbg_din_15_ ),
    .Y(_00671_)
  );
  OR2X1 _06496_ (
    .A( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .Y(_00672_)
  );
  AND2X1 _06497_ (
    .A( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .Y(_00673_)
  );
  OAI21X1 _06498_ (
    .A( dbg_0.dbg_i2c_0.scl_sync ),
    .B(_00673_),
    .C(_00672_),
    .Y(_00674_)
  );
  INVX1 _06499_ (
    .A(_00674_),
    .Y( dbg_0.dbg_i2c_0.scl )
  );
  OR2X1 _06500_ (
    .A( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .Y(_00675_)
  );
  AND2X1 _06501_ (
    .A( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .B( dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .Y(_00676_)
  );
  OAI21X1 _06502_ (
    .A( dbg_0.dbg_i2c_0.sda_in_sync ),
    .B(_00676_),
    .C(_00675_),
    .Y(_00677_)
  );
  INVX1 _06503_ (
    .A(_00677_),
    .Y( dbg_0.dbg_i2c_0.sda_in )
  );
  NOR3X1 _06504_ (
    .A(_00650_),
    .B(_00674_),
    .C( dbg_0.dbg_i2c_0.sda_in ),
    .Y(_00678_)
  );
  NAND3X1 _06505_ (
    .A( dbg_0.dbg_i2c_0.sda_in_dly ),
    .B( dbg_0.dbg_i2c_0.scl ),
    .C(_00677_),
    .Y(_00679_)
  );
  NOR3X1 _06506_ (
    .A( dbg_0.dbg_i2c_0.sda_in_dly ),
    .B(_00674_),
    .C(_00677_),
    .Y(_00680_)
  );
  NAND3X1 _06507_ (
    .A(_00650_),
    .B( dbg_0.dbg_i2c_0.scl ),
    .C( dbg_0.dbg_i2c_0.sda_in ),
    .Y(_00681_)
  );
  NOR2X1 _06508_ (
    .A(_00651_),
    .B(_00680_),
    .Y(_00682_)
  );
  NOR3X1 _06509_ (
    .A(_00651_),
    .B(_00678_),
    .C(_00680_),
    .Y(_00683_)
  );
  NAND3X1 _06510_ (
    .A( dbg_0.dbg_i2c_0.i2c_active_seq ),
    .B(_00679_),
    .C(_00681_),
    .Y(_00684_)
  );
  NOR2X1 _06511_ (
    .A(_00649_),
    .B( dbg_0.dbg_i2c_0.scl ),
    .Y(_00685_)
  );
  NAND2X1 _06512_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00674_),
    .Y(_00686_)
  );
  NOR3X1 _06513_ (
    .A(_00649_),
    .B(_00654_),
    .C( dbg_0.dbg_i2c_0.scl ),
    .Y(_00687_)
  );
  NAND3X1 _06514_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .C(_00674_),
    .Y(_00688_)
  );
  NOR2X1 _06515_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00689_)
  );
  NAND2X1 _06516_ (
    .A(_00652_),
    .B(_00653_),
    .Y(_00690_)
  );
  NAND3X1 _06517_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00687_),
    .C(_00689_),
    .Y(_00691_)
  );
  NOR2X1 _06518_ (
    .A(_00652_),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00692_)
  );
  OAI21X1 _06519_ (
    .A(_00677_),
    .B(_00688_),
    .C(_00692_),
    .Y(_00693_)
  );
  NAND2X1 _06520_ (
    .A(_00691_),
    .B(_00693_),
    .Y(_00694_)
  );
  AOI21X1 _06521_ (
    .A(_00691_),
    .B(_00693_),
    .C(_00684_),
    .Y( dbg_0.dbg_i2c_0.i2c_state_nxt_2_ )
  );
  NOR3X1 _06522_ (
    .A(_00649_),
    .B(_00656_),
    .C( dbg_0.dbg_i2c_0.scl ),
    .Y(_00695_)
  );
  NAND3X1 _06523_ (
    .A(_00654_),
    .B(_00689_),
    .C(_00695_),
    .Y(_00696_)
  );
  XOR2X1 _06524_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(dbg_i2c_addr_2_),
    .Y(_00697_)
  );
  NOR2X1 _06525_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_i2c_addr_5_),
    .Y(_00698_)
  );
  AND2X1 _06526_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_i2c_addr_5_),
    .Y(_00699_)
  );
  XNOR2X1 _06527_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(dbg_i2c_addr_4_),
    .Y(_00700_)
  );
  OAI21X1 _06528_ (
    .A(_00698_),
    .B(_00699_),
    .C(_00700_),
    .Y(_00701_)
  );
  NOR2X1 _06529_ (
    .A(_00697_),
    .B(_00701_),
    .Y(_00702_)
  );
  OAI22X1 _06530_ (
    .A(_00657_),
    .B(dbg_i2c_addr_0_),
    .C(dbg_i2c_addr_3_),
    .D(_00661_),
    .Y(_00703_)
  );
  XOR2X1 _06531_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(dbg_i2c_addr_6_),
    .Y(_00704_)
  );
  NOR2X1 _06532_ (
    .A(_00703_),
    .B(_00704_),
    .Y(_00705_)
  );
  XNOR2X1 _06533_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_i2c_addr_1_),
    .Y(_00706_)
  );
  AOI22X1 _06534_ (
    .A(_00657_),
    .B(dbg_i2c_addr_0_),
    .C(dbg_i2c_addr_3_),
    .D(_00661_),
    .Y(_00707_)
  );
  AND2X1 _06535_ (
    .A(_00706_),
    .B(_00707_),
    .Y(_00708_)
  );
  NAND3X1 _06536_ (
    .A(_00702_),
    .B(_00705_),
    .C(_00708_),
    .Y(_00709_)
  );
  INVX1 _06537_ (
    .A(_00709_),
    .Y(_00710_)
  );
  NAND2X1 _06538_ (
    .A(_00652_),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00711_)
  );
  OR2X1 _06539_ (
    .A(_00654_),
    .B(_00711_),
    .Y(_00712_)
  );
  AOI21X1 _06540_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .C(_00654_),
    .Y(_00713_)
  );
  NOR2X1 _06541_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .B(_00711_),
    .Y(_00714_)
  );
  AND2X1 _06542_ (
    .A(_00695_),
    .B(_00714_),
    .Y(_00715_)
  );
  NAND2X1 _06543_ (
    .A(_00695_),
    .B(_00714_),
    .Y(_00716_)
  );
  AOI22X1 _06544_ (
    .A(_00686_),
    .B(_00713_),
    .C(_00714_),
    .D(_00695_),
    .Y(_00717_)
  );
  OAI21X1 _06545_ (
    .A(_00696_),
    .B(_00709_),
    .C(_00717_),
    .Y(_00718_)
  );
  NOR2X1 _06546_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00719_)
  );
  NAND2X1 _06547_ (
    .A(_00655_),
    .B( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .Y(_00720_)
  );
  NOR2X1 _06548_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00721_)
  );
  NAND3X1 _06549_ (
    .A(_00657_),
    .B(_00658_),
    .C(_00721_),
    .Y(_00722_)
  );
  NOR2X1 _06550_ (
    .A(_00720_),
    .B(_00722_),
    .Y(_00723_)
  );
  NAND3X1 _06551_ (
    .A(_00663_),
    .B(_00719_),
    .C(_00723_),
    .Y(_00724_)
  );
  NAND2X1 _06552_ (
    .A(_00685_),
    .B(_00692_),
    .Y(_00725_)
  );
  NOR2X1 _06553_ (
    .A(_00724_),
    .B(_00725_),
    .Y(_00726_)
  );
  OR2X1 _06554_ (
    .A(_00724_),
    .B(_00725_),
    .Y(_00727_)
  );
  AOI21X1 _06555_ (
    .A(_00654_),
    .B(_00726_),
    .C(_00718_),
    .Y(_00728_)
  );
  NOR2X1 _06556_ (
    .A(_00684_),
    .B(_00728_),
    .Y( dbg_0.dbg_i2c_0.i2c_state_nxt_0_ )
  );
  NOR3X1 _06557_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00688_),
    .C(_00690_),
    .Y(_00729_)
  );
  NAND3X1 _06558_ (
    .A(_00655_),
    .B(_00687_),
    .C(_00689_),
    .Y(_00730_)
  );
  AOI21X1 _06559_ (
    .A(_00711_),
    .B(_00730_),
    .C(_00684_),
    .Y( dbg_0.dbg_i2c_0.i2c_state_nxt_1_ )
  );
  NOR2X1 _06560_ (
    .A( dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00674_),
    .Y( dbg_0.dbg_i2c_0.scl_re )
  );
  NOR2X1 _06561_ (
    .A(_00665_),
    .B(_00666_),
    .Y(_00731_)
  );
  AOI21X1 _06562_ (
    .A(_00665_),
    .B( dbg_0.dbg_i2c_0.dbg_bw ),
    .C(_00731_),
    .Y(_00732_)
  );
  NAND2X1 _06563_ (
    .A(_00664_),
    .B( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .Y(_00733_)
  );
  NOR2X1 _06564_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00733_),
    .Y(_00734_)
  );
  AND2X1 _06565_ (
    .A(_00715_),
    .B(_00734_),
    .Y(_00735_)
  );
  NOR2X1 _06566_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .Y(_00736_)
  );
  NAND2X1 _06567_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00736_),
    .Y(_00737_)
  );
  NOR2X1 _06568_ (
    .A(_00716_),
    .B(_00737_),
    .Y(_00738_)
  );
  MUX2X1 _06569_ (
    .A(_00735_),
    .B(_00738_),
    .S(_00732_),
    .Y(_00739_)
  );
  INVX1 _06570_ (
    .A(_00739_),
    .Y(_00613_)
  );
  NOR2X1 _06571_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .Y(_00740_)
  );
  AND2X1 _06572_ (
    .A(_00664_),
    .B(_00740_),
    .Y(_00741_)
  );
  AND2X1 _06573_ (
    .A(_00715_),
    .B(_00741_),
    .Y(_00742_)
  );
  NAND2X1 _06574_ (
    .A(_00715_),
    .B(_00741_),
    .Y(_00743_)
  );
  NAND2X1 _06575_ (
    .A(_00662_),
    .B(_00742_),
    .Y(_00744_)
  );
  NAND2X1 _06576_ (
    .A( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B(_00740_),
    .Y(_00745_)
  );
  NOR2X1 _06577_ (
    .A(_00665_),
    .B(_00745_),
    .Y(_00746_)
  );
  AND2X1 _06578_ (
    .A(_00726_),
    .B(_00746_),
    .Y(_00747_)
  );
  NAND3X1 _06579_ (
    .A(_00664_),
    .B( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .C( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .Y(_00748_)
  );
  INVX1 _06580_ (
    .A(_00748_),
    .Y(_00749_)
  );
  NOR2X1 _06581_ (
    .A(_00727_),
    .B(_00748_),
    .Y(_00750_)
  );
  AOI22X1 _06582_ (
    .A(_00666_),
    .B(_00747_),
    .C(_00750_),
    .D(_00731_),
    .Y(_00751_)
  );
  OAI21X1 _06583_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00744_),
    .C(_00751_),
    .Y(_00612_)
  );
  OAI21X1 _06584_ (
    .A(_00665_),
    .B(_00666_),
    .C(_00726_),
    .Y(_00752_)
  );
  AOI21X1 _06585_ (
    .A(_00749_),
    .B(_00752_),
    .C(_00747_),
    .Y(_00753_)
  );
  OR2X1 _06586_ (
    .A(_00665_),
    .B( dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00754_)
  );
  INVX1 _06587_ (
    .A(_00754_),
    .Y(_00755_)
  );
  OAI21X1 _06588_ (
    .A(_00666_),
    .B(_00754_),
    .C(_00715_),
    .Y(_00756_)
  );
  AOI21X1 _06589_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B( dbg_0.dbg_i2c_0.mem_burst_end ),
    .C(_00737_),
    .Y(_00757_)
  );
  OR2X1 _06590_ (
    .A( dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B( dbg_0.dbg_i2c_0.mem_burst_wr ),
    .Y(_00758_)
  );
  OAI21X1 _06591_ (
    .A(_00715_),
    .B(_00758_),
    .C(_00741_),
    .Y(_00759_)
  );
  AOI22X1 _06592_ (
    .A(_00735_),
    .B(_00755_),
    .C(_00756_),
    .D(_00757_),
    .Y(_00760_)
  );
  NAND3X1 _06593_ (
    .A(_00753_),
    .B(_00759_),
    .C(_00760_),
    .Y( dbg_0.dbg_i2c_0.dbg_state_nxt_0_ )
  );
  AOI22X1 _06594_ (
    .A( dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B(_00741_),
    .C(_00742_),
    .D(_00662_),
    .Y(_00761_)
  );
  OR2X1 _06595_ (
    .A( dbg_0.dbg_i2c_0.mem_burst_wr ),
    .B(_00761_),
    .Y(_00762_)
  );
  AOI21X1 _06596_ (
    .A(_00665_),
    .B( dbg_0.dbg_i2c_0.dbg_bw ),
    .C(_00756_),
    .Y(_00763_)
  );
  AOI22X1 _06597_ (
    .A(_00716_),
    .B(_00734_),
    .C(_00757_),
    .D(_00763_),
    .Y(_00764_)
  );
  NAND3X1 _06598_ (
    .A(_00753_),
    .B(_00762_),
    .C(_00764_),
    .Y( dbg_0.dbg_i2c_0.dbg_state_nxt_1_ )
  );
  NAND2X1 _06599_ (
    .A(_00732_),
    .B(_00750_),
    .Y(_00765_)
  );
  OAI21X1 _06600_ (
    .A(_00726_),
    .B(_00745_),
    .C(_00765_),
    .Y( dbg_0.dbg_i2c_0.dbg_state_nxt_2_ )
  );
  MUX2X1 _06601_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B( dbg_0.dbg_din_8_ ),
    .S(_00735_),
    .Y(_00766_)
  );
  NOR2X1 _06602_ (
    .A(_00738_),
    .B(_00766_),
    .Y(_00615_)
  );
  MUX2X1 _06603_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B( dbg_0.dbg_din_9_ ),
    .S(_00735_),
    .Y(_00767_)
  );
  NOR2X1 _06604_ (
    .A(_00738_),
    .B(_00767_),
    .Y(_00616_)
  );
  MUX2X1 _06605_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B( dbg_0.dbg_din_10_ ),
    .S(_00735_),
    .Y(_00768_)
  );
  NOR2X1 _06606_ (
    .A(_00738_),
    .B(_00768_),
    .Y(_00617_)
  );
  OR2X1 _06607_ (
    .A(_00735_),
    .B(_00738_),
    .Y(_00769_)
  );
  NAND2X1 _06608_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00735_),
    .Y(_00770_)
  );
  OAI21X1 _06609_ (
    .A(_00667_),
    .B(_00769_),
    .C(_00770_),
    .Y(_00618_)
  );
  NAND2X1 _06610_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00735_),
    .Y(_00771_)
  );
  OAI21X1 _06611_ (
    .A(_00668_),
    .B(_00769_),
    .C(_00771_),
    .Y(_00619_)
  );
  NAND2X1 _06612_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00735_),
    .Y(_00772_)
  );
  OAI21X1 _06613_ (
    .A(_00669_),
    .B(_00769_),
    .C(_00772_),
    .Y(_00620_)
  );
  NAND2X1 _06614_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00735_),
    .Y(_00773_)
  );
  OAI21X1 _06615_ (
    .A(_00670_),
    .B(_00769_),
    .C(_00773_),
    .Y(_00621_)
  );
  NAND2X1 _06616_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00735_),
    .Y(_00774_)
  );
  OAI21X1 _06617_ (
    .A(_00671_),
    .B(_00769_),
    .C(_00774_),
    .Y(_00622_)
  );
  NAND2X1 _06618_ (
    .A(_00655_),
    .B(_00738_),
    .Y(_00775_)
  );
  OAI21X1 _06619_ (
    .A( dbg_0.dbg_din_0_ ),
    .B(_00738_),
    .C(_00775_),
    .Y(_00776_)
  );
  INVX1 _06620_ (
    .A(_00776_),
    .Y(_00623_)
  );
  NAND2X1 _06621_ (
    .A(_00657_),
    .B(_00738_),
    .Y(_00777_)
  );
  OAI21X1 _06622_ (
    .A( dbg_0.dbg_din_1_ ),
    .B(_00738_),
    .C(_00777_),
    .Y(_00778_)
  );
  INVX1 _06623_ (
    .A(_00778_),
    .Y(_00624_)
  );
  NAND2X1 _06624_ (
    .A(_00659_),
    .B(_00738_),
    .Y(_00779_)
  );
  OAI21X1 _06625_ (
    .A( dbg_0.dbg_din_2_ ),
    .B(_00738_),
    .C(_00779_),
    .Y(_00780_)
  );
  INVX1 _06626_ (
    .A(_00780_),
    .Y(_00625_)
  );
  NAND2X1 _06627_ (
    .A(_00658_),
    .B(_00738_),
    .Y(_00781_)
  );
  OAI21X1 _06628_ (
    .A( dbg_0.dbg_din_3_ ),
    .B(_00738_),
    .C(_00781_),
    .Y(_00782_)
  );
  INVX1 _06629_ (
    .A(_00782_),
    .Y(_00626_)
  );
  NAND2X1 _06630_ (
    .A(_00661_),
    .B(_00738_),
    .Y(_00783_)
  );
  OAI21X1 _06631_ (
    .A( dbg_0.dbg_din_4_ ),
    .B(_00738_),
    .C(_00783_),
    .Y(_00784_)
  );
  INVX1 _06632_ (
    .A(_00784_),
    .Y(_00627_)
  );
  NAND2X1 _06633_ (
    .A(_00660_),
    .B(_00738_),
    .Y(_00785_)
  );
  OAI21X1 _06634_ (
    .A( dbg_0.dbg_din_5_ ),
    .B(_00738_),
    .C(_00785_),
    .Y(_00786_)
  );
  INVX1 _06635_ (
    .A(_00786_),
    .Y(_00628_)
  );
  NAND2X1 _06636_ (
    .A(_00663_),
    .B(_00738_),
    .Y(_00787_)
  );
  OAI21X1 _06637_ (
    .A( dbg_0.dbg_din_6_ ),
    .B(_00738_),
    .C(_00787_),
    .Y(_00788_)
  );
  INVX1 _06638_ (
    .A(_00788_),
    .Y(_00629_)
  );
  NAND2X1 _06639_ (
    .A(_00662_),
    .B(_00738_),
    .Y(_00789_)
  );
  OAI21X1 _06640_ (
    .A( dbg_0.dbg_din_7_ ),
    .B(_00738_),
    .C(_00789_),
    .Y(_00790_)
  );
  INVX1 _06641_ (
    .A(_00790_),
    .Y(_00630_)
  );
  NOR2X1 _06642_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00742_),
    .Y(_00791_)
  );
  OR2X1 _06643_ (
    .A( dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00742_),
    .Y(_00792_)
  );
  AOI22X1 _06644_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00742_),
    .C(_00791_),
    .D( dbg_0.dbg_addr_0_ ),
    .Y(_00793_)
  );
  INVX1 _06645_ (
    .A(_00793_),
    .Y(_00631_)
  );
  OAI22X1 _06646_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(_00743_),
    .C(_00792_),
    .D( dbg_0.dbg_addr_1_ ),
    .Y(_00794_)
  );
  INVX1 _06647_ (
    .A(_00794_),
    .Y(_00632_)
  );
  OAI22X1 _06648_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(_00743_),
    .C(_00792_),
    .D( dbg_0.dbg_addr_2_ ),
    .Y(_00795_)
  );
  INVX1 _06649_ (
    .A(_00795_),
    .Y(_00633_)
  );
  AOI22X1 _06650_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00742_),
    .C(_00791_),
    .D( dbg_0.dbg_addr_3_ ),
    .Y(_00796_)
  );
  INVX1 _06651_ (
    .A(_00796_),
    .Y(_00634_)
  );
  AOI22X1 _06652_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00742_),
    .C(_00791_),
    .D( dbg_0.dbg_addr_4_ ),
    .Y(_00797_)
  );
  INVX1 _06653_ (
    .A(_00797_),
    .Y(_00635_)
  );
  AOI22X1 _06654_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00742_),
    .C(_00791_),
    .D( dbg_0.dbg_addr_5_ ),
    .Y(_00798_)
  );
  INVX1 _06655_ (
    .A(_00798_),
    .Y(_00636_)
  );
  NAND2X1 _06656_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00742_),
    .Y(_00799_)
  );
  OAI21X1 _06657_ (
    .A(_00732_),
    .B(_00742_),
    .C(_00799_),
    .Y(_00637_)
  );
  NAND3X1 _06658_ (
    .A(_00685_),
    .B( dbg_0.dbg_i2c_0.i2c_state_nxt_2_ ),
    .C(_00724_),
    .Y(_00800_)
  );
  OAI21X1 _06659_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .B(_00654_),
    .C( dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .Y(_00801_)
  );
  NOR2X1 _06660_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B(_00801_),
    .Y(_00802_)
  );
  NOR2X1 _06661_ (
    .A(_00686_),
    .B(_00712_),
    .Y(_00803_)
  );
  OR2X1 _06662_ (
    .A(_00686_),
    .B(_00712_),
    .Y(_00804_)
  );
  NOR3X1 _06663_ (
    .A(_00684_),
    .B(_00729_),
    .C(_00803_),
    .Y(_00805_)
  );
  NAND3X1 _06664_ (
    .A(_00683_),
    .B(_00730_),
    .C(_00804_),
    .Y(_00806_)
  );
  NOR2X1 _06665_ (
    .A( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .Y(_00807_)
  );
  NAND3X1 _06666_ (
    .A(_00653_),
    .B( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .C( dbg_0.dbg_i2c_0.scl_re ),
    .Y(_00808_)
  );
  NOR2X1 _06667_ (
    .A(_00807_),
    .B(_00808_),
    .Y(_00809_)
  );
  OR2X1 _06668_ (
    .A(_00807_),
    .B(_00808_),
    .Y(_00810_)
  );
  OAI21X1 _06669_ (
    .A(_00807_),
    .B(_00808_),
    .C(_00805_),
    .Y(_00811_)
  );
  NOR3X1 _06670_ (
    .A(_00802_),
    .B(_00806_),
    .C(_00809_),
    .Y(_00812_)
  );
  AND2X1 _06671_ (
    .A(_00800_),
    .B(_00812_),
    .Y(_00813_)
  );
  NAND3X1 _06672_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00800_),
    .C(_00812_),
    .Y(_00814_)
  );
  NOR2X1 _06673_ (
    .A( dbg_0.dbg_i2c_0.sda_in ),
    .B(_00811_),
    .Y(_00815_)
  );
  OAI21X1 _06674_ (
    .A(_00812_),
    .B(_00815_),
    .C(_00814_),
    .Y(_00639_)
  );
  NAND2X1 _06675_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00808_),
    .Y(_00816_)
  );
  MUX2X1 _06676_ (
    .A( dbg_0.dbg_dout_0_ ),
    .B( dbg_0.dbg_dout_8_ ),
    .S(_00745_),
    .Y(_00817_)
  );
  OAI21X1 _06677_ (
    .A(_00810_),
    .B(_00817_),
    .C(_00816_),
    .Y(_00818_)
  );
  NAND2X1 _06678_ (
    .A(_00805_),
    .B(_00818_),
    .Y(_00819_)
  );
  MUX2X1 _06679_ (
    .A(_00657_),
    .B(_00819_),
    .S(_00813_),
    .Y(_00640_)
  );
  MUX2X1 _06680_ (
    .A( dbg_0.dbg_dout_1_ ),
    .B( dbg_0.dbg_dout_9_ ),
    .S(_00745_),
    .Y(_00820_)
  );
  MUX2X1 _06681_ (
    .A(_00657_),
    .B(_00820_),
    .S(_00810_),
    .Y(_00821_)
  );
  NAND2X1 _06682_ (
    .A(_00805_),
    .B(_00821_),
    .Y(_00822_)
  );
  MUX2X1 _06683_ (
    .A(_00659_),
    .B(_00822_),
    .S(_00813_),
    .Y(_00641_)
  );
  MUX2X1 _06684_ (
    .A( dbg_0.dbg_dout_2_ ),
    .B( dbg_0.dbg_dout_10_ ),
    .S(_00745_),
    .Y(_00823_)
  );
  MUX2X1 _06685_ (
    .A(_00659_),
    .B(_00823_),
    .S(_00810_),
    .Y(_00824_)
  );
  NAND2X1 _06686_ (
    .A(_00805_),
    .B(_00824_),
    .Y(_00825_)
  );
  MUX2X1 _06687_ (
    .A(_00658_),
    .B(_00825_),
    .S(_00813_),
    .Y(_00642_)
  );
  MUX2X1 _06688_ (
    .A( dbg_0.dbg_dout_3_ ),
    .B( dbg_0.dbg_dout_11_ ),
    .S(_00745_),
    .Y(_00826_)
  );
  MUX2X1 _06689_ (
    .A(_00658_),
    .B(_00826_),
    .S(_00810_),
    .Y(_00827_)
  );
  NAND2X1 _06690_ (
    .A(_00805_),
    .B(_00827_),
    .Y(_00828_)
  );
  MUX2X1 _06691_ (
    .A(_00661_),
    .B(_00828_),
    .S(_00813_),
    .Y(_00643_)
  );
  MUX2X1 _06692_ (
    .A( dbg_0.dbg_dout_4_ ),
    .B( dbg_0.dbg_dout_12_ ),
    .S(_00745_),
    .Y(_00829_)
  );
  MUX2X1 _06693_ (
    .A(_00661_),
    .B(_00829_),
    .S(_00810_),
    .Y(_00830_)
  );
  NAND2X1 _06694_ (
    .A(_00805_),
    .B(_00830_),
    .Y(_00831_)
  );
  MUX2X1 _06695_ (
    .A(_00660_),
    .B(_00831_),
    .S(_00813_),
    .Y(_00644_)
  );
  MUX2X1 _06696_ (
    .A( dbg_0.dbg_dout_5_ ),
    .B( dbg_0.dbg_dout_13_ ),
    .S(_00745_),
    .Y(_00832_)
  );
  MUX2X1 _06697_ (
    .A(_00660_),
    .B(_00832_),
    .S(_00810_),
    .Y(_00833_)
  );
  NAND2X1 _06698_ (
    .A(_00805_),
    .B(_00833_),
    .Y(_00834_)
  );
  MUX2X1 _06699_ (
    .A(_00663_),
    .B(_00834_),
    .S(_00813_),
    .Y(_00645_)
  );
  MUX2X1 _06700_ (
    .A( dbg_0.dbg_dout_6_ ),
    .B( dbg_0.dbg_dout_14_ ),
    .S(_00745_),
    .Y(_00835_)
  );
  MUX2X1 _06701_ (
    .A(_00663_),
    .B(_00835_),
    .S(_00810_),
    .Y(_00836_)
  );
  NAND2X1 _06702_ (
    .A(_00805_),
    .B(_00836_),
    .Y(_00837_)
  );
  MUX2X1 _06703_ (
    .A(_00662_),
    .B(_00837_),
    .S(_00813_),
    .Y(_00646_)
  );
  MUX2X1 _06704_ (
    .A( dbg_0.dbg_dout_7_ ),
    .B( dbg_0.dbg_dout_15_ ),
    .S(_00745_),
    .Y(_00838_)
  );
  MUX2X1 _06705_ (
    .A(_00662_),
    .B(_00838_),
    .S(_00810_),
    .Y(_00839_)
  );
  NAND2X1 _06706_ (
    .A(_00805_),
    .B(_00839_),
    .Y(_00840_)
  );
  MUX2X1 _06707_ (
    .A(_00656_),
    .B(_00840_),
    .S(_00813_),
    .Y(_00647_)
  );
  OAI21X1 _06708_ (
    .A(_00696_),
    .B(_00710_),
    .C(_00682_),
    .Y(_00841_)
  );
  NAND2X1 _06709_ (
    .A(_00679_),
    .B(_00841_),
    .Y(_00648_)
  );
  NOR3X1 _06710_ (
    .A(_00684_),
    .B(_00694_),
    .C(_00728_),
    .Y(_00842_)
  );
  OAI21X1 _06711_ (
    .A( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00800_),
    .C(_00685_),
    .Y(_00843_)
  );
  OAI21X1 _06712_ (
    .A(_00649_),
    .B( dbg_0.dbg_i2c_0.scl ),
    .C(_05583_),
    .Y(_00844_)
  );
  OAI21X1 _06713_ (
    .A(_00842_),
    .B(_00843_),
    .C(_00844_),
    .Y(_00638_)
  );
  DFFSR _06714_ (
    .CLK(dco_clk),
    .D(_00612_),
    .Q( dbg_0.dbg_i2c_0.dbg_rd ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06715_ (
    .CLK(dco_clk),
    .D(_00613_),
    .Q( dbg_0.dbg_i2c_0.dbg_wr ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06716_ (
    .CLK(dco_clk),
    .D(_00615_),
    .Q( dbg_0.dbg_din_8_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06717_ (
    .CLK(dco_clk),
    .D(_00616_),
    .Q( dbg_0.dbg_din_9_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06718_ (
    .CLK(dco_clk),
    .D(_00617_),
    .Q( dbg_0.dbg_din_10_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06719_ (
    .CLK(dco_clk),
    .D(_00618_),
    .Q( dbg_0.dbg_din_11_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06720_ (
    .CLK(dco_clk),
    .D(_00619_),
    .Q( dbg_0.dbg_din_12_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06721_ (
    .CLK(dco_clk),
    .D(_00620_),
    .Q( dbg_0.dbg_din_13_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06722_ (
    .CLK(dco_clk),
    .D(_00621_),
    .Q( dbg_0.dbg_din_14_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06723_ (
    .CLK(dco_clk),
    .D(_00622_),
    .Q( dbg_0.dbg_din_15_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06724_ (
    .CLK(dco_clk),
    .D(_00623_),
    .Q( dbg_0.dbg_din_0_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06725_ (
    .CLK(dco_clk),
    .D(_00624_),
    .Q( dbg_0.dbg_din_1_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06726_ (
    .CLK(dco_clk),
    .D(_00625_),
    .Q( dbg_0.dbg_din_2_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06727_ (
    .CLK(dco_clk),
    .D(_00626_),
    .Q( dbg_0.dbg_din_3_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06728_ (
    .CLK(dco_clk),
    .D(_00627_),
    .Q( dbg_0.dbg_din_4_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06729_ (
    .CLK(dco_clk),
    .D(_00628_),
    .Q( dbg_0.dbg_din_5_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06730_ (
    .CLK(dco_clk),
    .D(_00629_),
    .Q( dbg_0.dbg_din_6_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06731_ (
    .CLK(dco_clk),
    .D(_00630_),
    .Q( dbg_0.dbg_din_7_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06732_ (
    .CLK(dco_clk),
    .D(_00631_),
    .Q( dbg_0.dbg_addr_0_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06733_ (
    .CLK(dco_clk),
    .D(_00632_),
    .Q( dbg_0.dbg_addr_1_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06734_ (
    .CLK(dco_clk),
    .D(_00633_),
    .Q( dbg_0.dbg_addr_2_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06735_ (
    .CLK(dco_clk),
    .D(_00634_),
    .Q( dbg_0.dbg_addr_3_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06736_ (
    .CLK(dco_clk),
    .D(_00635_),
    .Q( dbg_0.dbg_addr_4_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06737_ (
    .CLK(dco_clk),
    .D(_00636_),
    .Q( dbg_0.dbg_addr_5_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06738_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.dbg_state_nxt_0_ ),
    .Q( dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06739_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.dbg_state_nxt_1_ ),
    .Q( dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06740_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.dbg_state_nxt_2_ ),
    .Q( dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06741_ (
    .CLK(dco_clk),
    .D(_00637_),
    .Q( dbg_0.dbg_i2c_0.dbg_bw ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06742_ (
    .CLK(dco_clk),
    .D(_00638_),
    .Q(_05583_),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06743_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.i2c_state_nxt_0_ ),
    .Q( dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06744_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.i2c_state_nxt_1_ ),
    .Q( dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06745_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.i2c_state_nxt_2_ ),
    .Q( dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06746_ (
    .CLK(dco_clk),
    .D(_00639_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06747_ (
    .CLK(dco_clk),
    .D(_00640_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06748_ (
    .CLK(dco_clk),
    .D(_00641_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06749_ (
    .CLK(dco_clk),
    .D(_00642_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06750_ (
    .CLK(dco_clk),
    .D(_00643_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06751_ (
    .CLK(dco_clk),
    .D(_00644_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06752_ (
    .CLK(dco_clk),
    .D(_00645_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06753_ (
    .CLK(dco_clk),
    .D(_00646_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06754_ (
    .CLK(dco_clk),
    .D(_00647_),
    .Q( dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06755_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_re ),
    .Q( dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06756_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .Q( dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .R(_00614_),
    .S(1'h1)
  );
  DFFSR _06757_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl ),
    .Q( dbg_0.dbg_i2c_0.scl_dly ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06758_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sda_in ),
    .Q( dbg_0.dbg_i2c_0.sda_in_dly ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06759_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sda_in_sync ),
    .Q( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06760_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Q( dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06761_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_sync ),
    .Q( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06762_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Q( dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .R(1'h1),
    .S(_00614_)
  );
  DFFSR _06763_ (
    .CLK(dco_clk),
    .D(_00648_),
    .Q( dbg_0.dbg_i2c_0.i2c_active_seq ),
    .R(_00614_),
    .S(1'h1)
  );
  INVX1 _06764_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00845_)
  );
  DFFSR _06765_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ),
    .Q( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .R(_00845_),
    .S(1'h1)
  );
  DFFSR _06766_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .Q( dbg_0.dbg_i2c_0.scl_sync_n ),
    .R(_00845_),
    .S(1'h1)
  );
  INVX1 _06767_ (
    .A( clock_module_0.dbg_rst ),
    .Y(_00846_)
  );
  DFFSR _06768_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ),
    .Q( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .R(_00846_),
    .S(1'h1)
  );
  DFFSR _06769_ (
    .CLK(dco_clk),
    .D( dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .Q( dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .R(_00846_),
    .S(1'h1)
  );
  INVX1 _06770_ (
    .A( execution_unit_0.e_state_0_ ),
    .Y(_00883_)
  );
  INVX1 _06771_ (
    .A( execution_unit_0.e_state_2_ ),
    .Y(_00884_)
  );
  INVX1 _06772_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .Y(_00885_)
  );
  INVX1 _06773_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_00886_)
  );
  INVX1 _06774_ (
    .A( execution_unit_0.inst_as_1_ ),
    .Y(_00887_)
  );
  INVX1 _06775_ (
    .A( execution_unit_0.mdb_in_8_ ),
    .Y(_00888_)
  );
  INVX1 _06776_ (
    .A( execution_unit_0.mab_lsb ),
    .Y(_00889_)
  );
  INVX1 _06777_ (
    .A( execution_unit_0.mdb_in_9_ ),
    .Y(_00890_)
  );
  INVX1 _06778_ (
    .A( execution_unit_0.mdb_in_10_ ),
    .Y(_00891_)
  );
  INVX1 _06779_ (
    .A( execution_unit_0.mdb_in_11_ ),
    .Y(_00892_)
  );
  INVX1 _06780_ (
    .A( execution_unit_0.mdb_in_12_ ),
    .Y(_00893_)
  );
  INVX1 _06781_ (
    .A( execution_unit_0.mdb_in_13_ ),
    .Y(_00894_)
  );
  INVX1 _06782_ (
    .A( execution_unit_0.mdb_in_14_ ),
    .Y(_00895_)
  );
  INVX1 _06783_ (
    .A( execution_unit_0.mdb_in_15_ ),
    .Y(_00896_)
  );
  INVX1 _06784_ (
    .A( execution_unit_0.mdb_in_buf_8_ ),
    .Y(_00897_)
  );
  INVX1 _06785_ (
    .A( execution_unit_0.mdb_in_buf_9_ ),
    .Y(_00898_)
  );
  INVX1 _06786_ (
    .A( execution_unit_0.mdb_in_buf_10_ ),
    .Y(_00899_)
  );
  INVX1 _06787_ (
    .A( execution_unit_0.mdb_in_buf_11_ ),
    .Y(_00900_)
  );
  INVX1 _06788_ (
    .A( execution_unit_0.mdb_in_buf_12_ ),
    .Y(_00901_)
  );
  INVX1 _06789_ (
    .A( execution_unit_0.mdb_in_buf_13_ ),
    .Y(_00902_)
  );
  INVX1 _06790_ (
    .A( execution_unit_0.mdb_in_buf_14_ ),
    .Y(_00903_)
  );
  INVX1 _06791_ (
    .A( execution_unit_0.mdb_in_buf_15_ ),
    .Y(_00904_)
  );
  INVX1 _06792_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_00905_)
  );
  INVX1 _06793_ (
    .A( execution_unit_0.mdb_out_nxt_8_ ),
    .Y(_00906_)
  );
  INVX1 _06794_ (
    .A( execution_unit_0.mdb_out_nxt_9_ ),
    .Y(_00907_)
  );
  INVX1 _06795_ (
    .A( execution_unit_0.mdb_out_nxt_10_ ),
    .Y(_00908_)
  );
  INVX1 _06796_ (
    .A( execution_unit_0.mdb_out_nxt_11_ ),
    .Y(_00909_)
  );
  INVX1 _06797_ (
    .A( execution_unit_0.mdb_out_nxt_12_ ),
    .Y(_00910_)
  );
  INVX1 _06798_ (
    .A( execution_unit_0.mdb_out_nxt_13_ ),
    .Y(_00911_)
  );
  INVX1 _06799_ (
    .A( execution_unit_0.mdb_out_nxt_14_ ),
    .Y(_00912_)
  );
  INVX1 _06800_ (
    .A( execution_unit_0.mdb_out_nxt_15_ ),
    .Y(_00913_)
  );
  INVX1 _06801_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .Y(_00914_)
  );
  INVX1 _06802_ (
    .A( dbg_0.dbg_reg_wr ),
    .Y(_00915_)
  );
  INVX1 _06803_ (
    .A( execution_unit_0.inst_irq_rst ),
    .Y(_00916_)
  );
  INVX1 _06804_ (
    .A( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_00917_)
  );
  INVX1 _06805_ (
    .A(_05695_),
    .Y(_00848_)
  );
  AND2X1 _06806_ (
    .A(_00884_),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_00918_)
  );
  AND2X1 _06807_ (
    .A( execution_unit_0.e_state_1_ ),
    .B( execution_unit_0.e_state_0_ ),
    .Y(_00919_)
  );
  NAND3X1 _06808_ (
    .A(_00884_),
    .B( execution_unit_0.e_state_3_ ),
    .C(_00919_),
    .Y(_00920_)
  );
  INVX1 _06809_ (
    .A(_00920_),
    .Y( execution_unit_0.alu_0.exec_cycle )
  );
  NOR2X1 _06810_ (
    .A( execution_unit_0.e_state_2_ ),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_00921_)
  );
  NAND2X1 _06811_ (
    .A(_00883_),
    .B(_00921_),
    .Y(_00922_)
  );
  NOR2X1 _06812_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_00922_),
    .Y( execution_unit_0.reg_sr_clr )
  );
  NOR2X1 _06813_ (
    .A(_00884_),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_00923_)
  );
  NAND2X1 _06814_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_00923_),
    .Y(_00924_)
  );
  AND2X1 _06815_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_00883_),
    .Y(_00925_)
  );
  NAND2X1 _06816_ (
    .A(_00923_),
    .B(_00925_),
    .Y(_00926_)
  );
  INVX1 _06817_ (
    .A(_00926_),
    .Y(_00847_)
  );
  NOR2X1 _06818_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_00883_),
    .Y(_00927_)
  );
  AND2X1 _06819_ (
    .A(_00918_),
    .B(_00927_),
    .Y(_00928_)
  );
  NAND2X1 _06820_ (
    .A(_00918_),
    .B(_00927_),
    .Y(_00929_)
  );
  NOR2X1 _06821_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_00930_)
  );
  OR2X1 _06822_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_00931_)
  );
  NOR3X1 _06823_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_00883_),
    .C(_00930_),
    .Y(_00932_)
  );
  NAND2X1 _06824_ (
    .A(_00918_),
    .B(_00932_),
    .Y(_00933_)
  );
  NAND3X1 _06825_ (
    .A( execution_unit_0.inst_as_1_ ),
    .B(_00923_),
    .C(_00932_),
    .Y(_00934_)
  );
  OAI21X1 _06826_ (
    .A(_00929_),
    .B(_00930_),
    .C(_00934_),
    .Y(_00935_)
  );
  AOI21X1 _06827_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_00921_),
    .C(_00935_),
    .Y(_00936_)
  );
  NOR2X1 _06828_ (
    .A(_00886_),
    .B(_00929_),
    .Y( execution_unit_0.reg_sr_wr )
  );
  NOR2X1 _06829_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B( execution_unit_0.inst_as_2_ ),
    .Y(_00937_)
  );
  OR2X1 _06830_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B( execution_unit_0.inst_as_1_ ),
    .Y(_00938_)
  );
  NOR2X1 _06831_ (
    .A( execution_unit_0.inst_as_4_ ),
    .B(_00938_),
    .Y(_00939_)
  );
  AOI21X1 _06832_ (
    .A(_00937_),
    .B(_00939_),
    .C(_00920_),
    .Y(_00940_)
  );
  NOR2X1 _06833_ (
    .A( execution_unit_0.reg_sr_wr ),
    .B(_00940_),
    .Y(_00941_)
  );
  NAND2X1 _06834_ (
    .A(_00918_),
    .B(_00925_),
    .Y(_00942_)
  );
  NAND3X1 _06835_ (
    .A(_00886_),
    .B(_00918_),
    .C(_00925_),
    .Y(_00943_)
  );
  AOI21X1 _06836_ (
    .A(_00929_),
    .B(_00943_),
    .C(_00931_),
    .Y(_00944_)
  );
  NOR2X1 _06837_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( execution_unit_0.inst_as_7_ ),
    .Y(_00945_)
  );
  NOR2X1 _06838_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B( execution_unit_0.inst_as_5_ ),
    .Y(_00946_)
  );
  AOI21X1 _06839_ (
    .A(_00945_),
    .B(_00946_),
    .C(_00920_),
    .Y(_00947_)
  );
  AOI22X1 _06840_ (
    .A( execution_unit_0.inst_dext_0_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_0_ ),
    .Y(_00948_)
  );
  NAND2X1 _06841_ (
    .A( execution_unit_0.mab_lsb ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_00949_)
  );
  MUX2X1 _06842_ (
    .A( execution_unit_0.mdb_in_0_ ),
    .B( execution_unit_0.mdb_in_8_ ),
    .S(_00949_),
    .Y(_00950_)
  );
  NOR2X1 _06843_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00950_),
    .Y(_00951_)
  );
  AOI21X1 _06844_ (
    .A( execution_unit_0.mdb_in_buf_0_ ),
    .B( execution_unit_0.mdb_in_buf_valid ),
    .C(_00951_),
    .Y(_00952_)
  );
  MUX2X1 _06845_ (
    .A(_00948_),
    .B(_00952_),
    .S(_00941_),
    .Y(_00953_)
  );
  NOR2X1 _06846_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_00920_),
    .Y(_00954_)
  );
  AND2X1 _06847_ (
    .A( execution_unit_0.inst_as_0_ ),
    .B(_00954_),
    .Y(_00955_)
  );
  OAI21X1 _06848_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B(_00924_),
    .C(_00922_),
    .Y(_00956_)
  );
  OR2X1 _06849_ (
    .A(_00955_),
    .B(_00956_),
    .Y(_00957_)
  );
  MUX2X1 _06850_ (
    .A(_00953_),
    .B( dbg_0.dbg_reg_din_0_ ),
    .S(_00936_),
    .Y(_00958_)
  );
  OAI21X1 _06851_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_0_ ),
    .Y(_00959_)
  );
  OAI21X1 _06852_ (
    .A(_00957_),
    .B(_00958_),
    .C(_00959_),
    .Y( execution_unit_0.alu_0.alu_swpb_8_ )
  );
  AOI22X1 _06853_ (
    .A( execution_unit_0.inst_dext_1_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_1_ ),
    .Y(_00960_)
  );
  MUX2X1 _06854_ (
    .A( execution_unit_0.mdb_in_1_ ),
    .B( execution_unit_0.mdb_in_9_ ),
    .S(_00949_),
    .Y(_00961_)
  );
  NOR2X1 _06855_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00961_),
    .Y(_00962_)
  );
  AOI21X1 _06856_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_1_ ),
    .C(_00962_),
    .Y(_00963_)
  );
  MUX2X1 _06857_ (
    .A(_00960_),
    .B(_00963_),
    .S(_00941_),
    .Y(_00964_)
  );
  MUX2X1 _06858_ (
    .A(_00964_),
    .B( dbg_0.dbg_reg_din_1_ ),
    .S(_00936_),
    .Y(_00965_)
  );
  OAI21X1 _06859_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_1_ ),
    .Y(_00966_)
  );
  OAI21X1 _06860_ (
    .A(_00957_),
    .B(_00965_),
    .C(_00966_),
    .Y( execution_unit_0.alu_0.alu_shift_0_ )
  );
  AOI22X1 _06861_ (
    .A( execution_unit_0.inst_dext_2_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_2_ ),
    .Y(_00967_)
  );
  MUX2X1 _06862_ (
    .A( execution_unit_0.mdb_in_2_ ),
    .B( execution_unit_0.mdb_in_10_ ),
    .S(_00949_),
    .Y(_00968_)
  );
  NOR2X1 _06863_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00968_),
    .Y(_00969_)
  );
  AOI21X1 _06864_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_2_ ),
    .C(_00969_),
    .Y(_00970_)
  );
  MUX2X1 _06865_ (
    .A(_00967_),
    .B(_00970_),
    .S(_00941_),
    .Y(_00971_)
  );
  MUX2X1 _06866_ (
    .A(_00971_),
    .B( dbg_0.dbg_reg_din_2_ ),
    .S(_00936_),
    .Y(_00972_)
  );
  OAI21X1 _06867_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_2_ ),
    .Y(_00973_)
  );
  OAI21X1 _06868_ (
    .A(_00957_),
    .B(_00972_),
    .C(_00973_),
    .Y( execution_unit_0.alu_0.alu_shift_1_ )
  );
  AOI22X1 _06869_ (
    .A( execution_unit_0.inst_dext_3_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_3_ ),
    .Y(_00974_)
  );
  MUX2X1 _06870_ (
    .A( execution_unit_0.mdb_in_3_ ),
    .B( execution_unit_0.mdb_in_11_ ),
    .S(_00949_),
    .Y(_00975_)
  );
  NOR2X1 _06871_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00975_),
    .Y(_00976_)
  );
  AOI21X1 _06872_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_3_ ),
    .C(_00976_),
    .Y(_00977_)
  );
  MUX2X1 _06873_ (
    .A(_00974_),
    .B(_00977_),
    .S(_00941_),
    .Y(_00978_)
  );
  MUX2X1 _06874_ (
    .A(_00978_),
    .B( dbg_0.dbg_reg_din_3_ ),
    .S(_00936_),
    .Y(_00979_)
  );
  OAI21X1 _06875_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_3_ ),
    .Y(_00980_)
  );
  OAI21X1 _06876_ (
    .A(_00957_),
    .B(_00979_),
    .C(_00980_),
    .Y( execution_unit_0.alu_0.alu_shift_2_ )
  );
  AOI22X1 _06877_ (
    .A( execution_unit_0.inst_dext_4_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_4_ ),
    .Y(_00981_)
  );
  MUX2X1 _06878_ (
    .A( execution_unit_0.mdb_in_4_ ),
    .B( execution_unit_0.mdb_in_12_ ),
    .S(_00949_),
    .Y(_00982_)
  );
  NOR2X1 _06879_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00982_),
    .Y(_00983_)
  );
  AOI21X1 _06880_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_4_ ),
    .C(_00983_),
    .Y(_00984_)
  );
  MUX2X1 _06881_ (
    .A(_00981_),
    .B(_00984_),
    .S(_00941_),
    .Y(_00985_)
  );
  MUX2X1 _06882_ (
    .A(_00985_),
    .B( dbg_0.dbg_reg_din_4_ ),
    .S(_00936_),
    .Y(_00986_)
  );
  OAI21X1 _06883_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_4_ ),
    .Y(_00987_)
  );
  OAI21X1 _06884_ (
    .A(_00957_),
    .B(_00986_),
    .C(_00987_),
    .Y( execution_unit_0.alu_0.alu_shift_3_ )
  );
  AOI22X1 _06885_ (
    .A( execution_unit_0.inst_dext_5_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_5_ ),
    .Y(_00988_)
  );
  MUX2X1 _06886_ (
    .A( execution_unit_0.mdb_in_5_ ),
    .B( execution_unit_0.mdb_in_13_ ),
    .S(_00949_),
    .Y(_00989_)
  );
  NOR2X1 _06887_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00989_),
    .Y(_00990_)
  );
  AOI21X1 _06888_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_5_ ),
    .C(_00990_),
    .Y(_00991_)
  );
  MUX2X1 _06889_ (
    .A(_00988_),
    .B(_00991_),
    .S(_00941_),
    .Y(_00992_)
  );
  MUX2X1 _06890_ (
    .A(_00992_),
    .B( dbg_0.dbg_reg_din_5_ ),
    .S(_00936_),
    .Y(_00993_)
  );
  OAI21X1 _06891_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_5_ ),
    .Y(_00994_)
  );
  OAI21X1 _06892_ (
    .A(_00957_),
    .B(_00993_),
    .C(_00994_),
    .Y( execution_unit_0.alu_0.alu_shift_4_ )
  );
  AOI22X1 _06893_ (
    .A( execution_unit_0.inst_dext_6_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_6_ ),
    .Y(_00995_)
  );
  MUX2X1 _06894_ (
    .A( execution_unit_0.mdb_in_6_ ),
    .B( execution_unit_0.mdb_in_14_ ),
    .S(_00949_),
    .Y(_00996_)
  );
  NOR2X1 _06895_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_00996_),
    .Y(_00997_)
  );
  AOI21X1 _06896_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_6_ ),
    .C(_00997_),
    .Y(_00998_)
  );
  MUX2X1 _06897_ (
    .A(_00995_),
    .B(_00998_),
    .S(_00941_),
    .Y(_00999_)
  );
  MUX2X1 _06898_ (
    .A(_00999_),
    .B( dbg_0.dbg_reg_din_6_ ),
    .S(_00936_),
    .Y(_01000_)
  );
  OAI21X1 _06899_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_6_ ),
    .Y(_01001_)
  );
  OAI21X1 _06900_ (
    .A(_00957_),
    .B(_01000_),
    .C(_01001_),
    .Y( execution_unit_0.alu_0.alu_shift_5_ )
  );
  AOI22X1 _06901_ (
    .A( execution_unit_0.inst_dext_7_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_7_ ),
    .Y(_01002_)
  );
  MUX2X1 _06902_ (
    .A( execution_unit_0.mdb_in_7_ ),
    .B( execution_unit_0.mdb_in_15_ ),
    .S(_00949_),
    .Y(_01003_)
  );
  NOR2X1 _06903_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B(_01003_),
    .Y(_01004_)
  );
  AOI21X1 _06904_ (
    .A( execution_unit_0.mdb_in_buf_valid ),
    .B( execution_unit_0.mdb_in_buf_7_ ),
    .C(_01004_),
    .Y(_01005_)
  );
  MUX2X1 _06905_ (
    .A(_01002_),
    .B(_01005_),
    .S(_00941_),
    .Y(_01006_)
  );
  MUX2X1 _06906_ (
    .A(_01006_),
    .B( dbg_0.dbg_reg_din_7_ ),
    .S(_00936_),
    .Y(_01007_)
  );
  OAI21X1 _06907_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_7_ ),
    .Y(_01008_)
  );
  OAI21X1 _06908_ (
    .A(_00957_),
    .B(_01007_),
    .C(_01008_),
    .Y( execution_unit_0.alu_0.alu_shift_6_ )
  );
  AOI22X1 _06909_ (
    .A( execution_unit_0.inst_dext_8_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_8_ ),
    .Y(_01009_)
  );
  MUX2X1 _06910_ (
    .A( execution_unit_0.mdb_in_buf_8_ ),
    .B( execution_unit_0.mdb_in_8_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01010_)
  );
  MUX2X1 _06911_ (
    .A(_01009_),
    .B(_01010_),
    .S(_00941_),
    .Y(_01011_)
  );
  MUX2X1 _06912_ (
    .A(_01011_),
    .B( dbg_0.dbg_reg_din_8_ ),
    .S(_00936_),
    .Y(_01012_)
  );
  OAI21X1 _06913_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_8_ ),
    .Y(_01013_)
  );
  OAI21X1 _06914_ (
    .A(_00957_),
    .B(_01012_),
    .C(_01013_),
    .Y( execution_unit_0.alu_0.alu_swpb_0_ )
  );
  AOI22X1 _06915_ (
    .A( execution_unit_0.inst_dext_9_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_9_ ),
    .Y(_01014_)
  );
  MUX2X1 _06916_ (
    .A( execution_unit_0.mdb_in_buf_9_ ),
    .B( execution_unit_0.mdb_in_9_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01015_)
  );
  MUX2X1 _06917_ (
    .A(_01014_),
    .B(_01015_),
    .S(_00941_),
    .Y(_01016_)
  );
  MUX2X1 _06918_ (
    .A(_01016_),
    .B( dbg_0.dbg_reg_din_9_ ),
    .S(_00936_),
    .Y(_01017_)
  );
  OAI21X1 _06919_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_9_ ),
    .Y(_01018_)
  );
  OAI21X1 _06920_ (
    .A(_00957_),
    .B(_01017_),
    .C(_01018_),
    .Y( execution_unit_0.alu_0.alu_shift_8_ )
  );
  AOI22X1 _06921_ (
    .A( execution_unit_0.inst_dext_10_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_10_ ),
    .Y(_01019_)
  );
  MUX2X1 _06922_ (
    .A( execution_unit_0.mdb_in_buf_10_ ),
    .B( execution_unit_0.mdb_in_10_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01020_)
  );
  MUX2X1 _06923_ (
    .A(_01019_),
    .B(_01020_),
    .S(_00941_),
    .Y(_01021_)
  );
  MUX2X1 _06924_ (
    .A(_01021_),
    .B( dbg_0.dbg_reg_din_10_ ),
    .S(_00936_),
    .Y(_01022_)
  );
  OAI21X1 _06925_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_10_ ),
    .Y(_01023_)
  );
  OAI21X1 _06926_ (
    .A(_00957_),
    .B(_01022_),
    .C(_01023_),
    .Y( execution_unit_0.alu_0.alu_shift_9_ )
  );
  AOI22X1 _06927_ (
    .A( execution_unit_0.inst_dext_11_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_11_ ),
    .Y(_01024_)
  );
  MUX2X1 _06928_ (
    .A( execution_unit_0.mdb_in_buf_11_ ),
    .B( execution_unit_0.mdb_in_11_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01025_)
  );
  MUX2X1 _06929_ (
    .A(_01024_),
    .B(_01025_),
    .S(_00941_),
    .Y(_01026_)
  );
  MUX2X1 _06930_ (
    .A(_01026_),
    .B( dbg_0.dbg_reg_din_11_ ),
    .S(_00936_),
    .Y(_01027_)
  );
  OAI21X1 _06931_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_11_ ),
    .Y(_01028_)
  );
  OAI21X1 _06932_ (
    .A(_00957_),
    .B(_01027_),
    .C(_01028_),
    .Y( execution_unit_0.alu_0.alu_shift_10_ )
  );
  AOI22X1 _06933_ (
    .A( execution_unit_0.inst_dext_12_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_12_ ),
    .Y(_01029_)
  );
  MUX2X1 _06934_ (
    .A( execution_unit_0.mdb_in_buf_12_ ),
    .B( execution_unit_0.mdb_in_12_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01030_)
  );
  MUX2X1 _06935_ (
    .A(_01029_),
    .B(_01030_),
    .S(_00941_),
    .Y(_01031_)
  );
  MUX2X1 _06936_ (
    .A(_01031_),
    .B( dbg_0.dbg_reg_din_12_ ),
    .S(_00936_),
    .Y(_01032_)
  );
  OAI21X1 _06937_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_12_ ),
    .Y(_01033_)
  );
  OAI21X1 _06938_ (
    .A(_00957_),
    .B(_01032_),
    .C(_01033_),
    .Y( execution_unit_0.alu_0.alu_shift_11_ )
  );
  AOI22X1 _06939_ (
    .A( execution_unit_0.inst_dext_13_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_13_ ),
    .Y(_01034_)
  );
  MUX2X1 _06940_ (
    .A( execution_unit_0.mdb_in_buf_13_ ),
    .B( execution_unit_0.mdb_in_13_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01035_)
  );
  MUX2X1 _06941_ (
    .A(_01034_),
    .B(_01035_),
    .S(_00941_),
    .Y(_01036_)
  );
  MUX2X1 _06942_ (
    .A(_01036_),
    .B( dbg_0.dbg_reg_din_13_ ),
    .S(_00936_),
    .Y(_01037_)
  );
  OAI21X1 _06943_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_13_ ),
    .Y(_01038_)
  );
  OAI21X1 _06944_ (
    .A(_00957_),
    .B(_01037_),
    .C(_01038_),
    .Y( execution_unit_0.alu_0.alu_shift_12_ )
  );
  AOI22X1 _06945_ (
    .A( execution_unit_0.inst_dext_14_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_14_ ),
    .Y(_01039_)
  );
  MUX2X1 _06946_ (
    .A( execution_unit_0.mdb_in_buf_14_ ),
    .B( execution_unit_0.mdb_in_14_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01040_)
  );
  MUX2X1 _06947_ (
    .A(_01039_),
    .B(_01040_),
    .S(_00941_),
    .Y(_01041_)
  );
  MUX2X1 _06948_ (
    .A(_01041_),
    .B( dbg_0.dbg_reg_din_14_ ),
    .S(_00936_),
    .Y(_01042_)
  );
  OAI21X1 _06949_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_14_ ),
    .Y(_01043_)
  );
  OAI21X1 _06950_ (
    .A(_00957_),
    .B(_01042_),
    .C(_01043_),
    .Y( execution_unit_0.alu_0.alu_shift_13_ )
  );
  AOI22X1 _06951_ (
    .A( execution_unit_0.inst_dext_15_ ),
    .B(_00944_),
    .C(_00947_),
    .D( execution_unit_0.inst_sext_15_ ),
    .Y(_01044_)
  );
  MUX2X1 _06952_ (
    .A( execution_unit_0.mdb_in_buf_15_ ),
    .B( execution_unit_0.mdb_in_15_ ),
    .S( execution_unit_0.mdb_in_buf_valid ),
    .Y(_01045_)
  );
  MUX2X1 _06953_ (
    .A(_01044_),
    .B(_01045_),
    .S(_00941_),
    .Y(_01046_)
  );
  MUX2X1 _06954_ (
    .A(_01046_),
    .B( dbg_0.dbg_reg_din_15_ ),
    .S(_00936_),
    .Y(_01047_)
  );
  OAI21X1 _06955_ (
    .A(_00955_),
    .B(_00956_),
    .C( execution_unit_0.reg_src_15_ ),
    .Y(_01048_)
  );
  OAI21X1 _06956_ (
    .A(_00957_),
    .B(_01047_),
    .C(_01048_),
    .Y( execution_unit_0.alu_0.alu_shift_14_ )
  );
  OR2X1 _06957_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( execution_unit_0.inst_ad_0_ ),
    .Y(_01049_)
  );
  NOR2X1 _06958_ (
    .A( execution_unit_0.inst_type_0_ ),
    .B(_01049_),
    .Y(_01050_)
  );
  INVX1 _06959_ (
    .A(_01050_),
    .Y(_01051_)
  );
  OR2X1 _06960_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_00920_),
    .Y(_01052_)
  );
  NOR2X1 _06961_ (
    .A(_01050_),
    .B(_01052_),
    .Y(_01053_)
  );
  NOR2X1 _06962_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_00931_),
    .Y(_01054_)
  );
  NAND3X1 _06963_ (
    .A(_00918_),
    .B(_00927_),
    .C(_01054_),
    .Y(_01055_)
  );
  AOI21X1 _06964_ (
    .A(_00942_),
    .B(_01055_),
    .C( execution_unit_0.inst_ad_6_ ),
    .Y(_01056_)
  );
  NOR2X1 _06965_ (
    .A(_01053_),
    .B(_01056_),
    .Y(_01057_)
  );
  NOR2X1 _06966_ (
    .A(_01051_),
    .B(_01052_),
    .Y(_01058_)
  );
  NAND3X1 _06967_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_00918_),
    .C(_00925_),
    .Y(_01059_)
  );
  INVX1 _06968_ (
    .A(_01059_),
    .Y(_01060_)
  );
  NOR2X1 _06969_ (
    .A(_01058_),
    .B(_01060_),
    .Y(_01061_)
  );
  OAI21X1 _06970_ (
    .A(_01051_),
    .B(_01052_),
    .C(_01059_),
    .Y(_01062_)
  );
  NOR2X1 _06971_ (
    .A(_01057_),
    .B(_01062_),
    .Y(_01063_)
  );
  NOR2X1 _06972_ (
    .A(_00924_),
    .B(_00939_),
    .Y(_01064_)
  );
  OR2X1 _06973_ (
    .A(_00924_),
    .B(_00939_),
    .Y(_01065_)
  );
  NAND2X1 _06974_ (
    .A( execution_unit_0.inst_sext_0_ ),
    .B(_01064_),
    .Y(_01066_)
  );
  OAI21X1 _06975_ (
    .A(_00950_),
    .B(_01061_),
    .C(_01066_),
    .Y(_01067_)
  );
  AOI21X1 _06976_ (
    .A( dbg_0.dbg_reg_din_0_ ),
    .B(_01063_),
    .C(_01067_),
    .Y(_01068_)
  );
  NAND2X1 _06977_ (
    .A(_05677_),
    .B( dbg_0.cpu_stat_full_0_ ),
    .Y(_01069_)
  );
  OAI21X1 _06978_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01068_),
    .C(_01069_),
    .Y( execution_unit_0.alu_0.op_dst_0_ )
  );
  NAND2X1 _06979_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05684_),
    .Y(_01070_)
  );
  OAI21X1 _06980_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_1_ ),
    .Y(_01071_)
  );
  OAI21X1 _06981_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B( execution_unit_0.inst_as_2_ ),
    .C( execution_unit_0.inst_src_1_ ),
    .Y(_01072_)
  );
  OR2X1 _06982_ (
    .A(_00930_),
    .B(_01072_),
    .Y(_01073_)
  );
  OAI21X1 _06983_ (
    .A(_00926_),
    .B(_01073_),
    .C(_00934_),
    .Y(_01074_)
  );
  OAI21X1 _06984_ (
    .A( execution_unit_0.e_state_1_ ),
    .B( execution_unit_0.e_state_0_ ),
    .C(_00921_),
    .Y(_01075_)
  );
  OAI21X1 _06985_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_00933_),
    .C(_01075_),
    .Y(_01076_)
  );
  NOR3X1 _06986_ (
    .A(_01062_),
    .B(_01074_),
    .C(_01076_),
    .Y(_01077_)
  );
  AOI22X1 _06987_ (
    .A(_00961_),
    .B(_01062_),
    .C(_01071_),
    .D(_01077_),
    .Y(_01078_)
  );
  MUX2X1 _06988_ (
    .A( execution_unit_0.inst_sext_1_ ),
    .B(_01078_),
    .S(_01064_),
    .Y(_01079_)
  );
  OAI21X1 _06989_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01079_),
    .C(_01070_),
    .Y( execution_unit_0.alu_0.op_dst_1_ )
  );
  NAND2X1 _06990_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05685_),
    .Y(_01080_)
  );
  OAI21X1 _06991_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_2_ ),
    .Y(_01081_)
  );
  AOI22X1 _06992_ (
    .A(_00968_),
    .B(_01062_),
    .C(_01077_),
    .D(_01081_),
    .Y(_01082_)
  );
  MUX2X1 _06993_ (
    .A( execution_unit_0.inst_sext_2_ ),
    .B(_01082_),
    .S(_01064_),
    .Y(_01083_)
  );
  OAI21X1 _06994_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01083_),
    .C(_01080_),
    .Y( execution_unit_0.alu_0.op_dst_2_ )
  );
  NAND2X1 _06995_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05686_),
    .Y(_01084_)
  );
  OAI21X1 _06996_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_3_ ),
    .Y(_01085_)
  );
  AOI22X1 _06997_ (
    .A(_00975_),
    .B(_01062_),
    .C(_01077_),
    .D(_01085_),
    .Y(_01086_)
  );
  MUX2X1 _06998_ (
    .A( execution_unit_0.inst_sext_3_ ),
    .B(_01086_),
    .S(_01064_),
    .Y(_01087_)
  );
  OAI21X1 _06999_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01087_),
    .C(_01084_),
    .Y( execution_unit_0.alu_0.op_dst_3_ )
  );
  NAND2X1 _07000_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05687_),
    .Y(_01088_)
  );
  OAI21X1 _07001_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_4_ ),
    .Y(_01089_)
  );
  AOI22X1 _07002_ (
    .A(_00982_),
    .B(_01062_),
    .C(_01077_),
    .D(_01089_),
    .Y(_01090_)
  );
  MUX2X1 _07003_ (
    .A( execution_unit_0.inst_sext_4_ ),
    .B(_01090_),
    .S(_01064_),
    .Y(_01091_)
  );
  OAI21X1 _07004_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01091_),
    .C(_01088_),
    .Y( execution_unit_0.alu_0.op_dst_4_ )
  );
  NAND2X1 _07005_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05688_),
    .Y(_01092_)
  );
  OAI21X1 _07006_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_5_ ),
    .Y(_01093_)
  );
  AOI22X1 _07007_ (
    .A(_00989_),
    .B(_01062_),
    .C(_01077_),
    .D(_01093_),
    .Y(_01094_)
  );
  MUX2X1 _07008_ (
    .A( execution_unit_0.inst_sext_5_ ),
    .B(_01094_),
    .S(_01064_),
    .Y(_01095_)
  );
  OAI21X1 _07009_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01095_),
    .C(_01092_),
    .Y( execution_unit_0.alu_0.op_dst_5_ )
  );
  NAND2X1 _07010_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05689_),
    .Y(_01096_)
  );
  OAI21X1 _07011_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_6_ ),
    .Y(_01097_)
  );
  AOI22X1 _07012_ (
    .A(_00996_),
    .B(_01062_),
    .C(_01077_),
    .D(_01097_),
    .Y(_01098_)
  );
  MUX2X1 _07013_ (
    .A( execution_unit_0.inst_sext_6_ ),
    .B(_01098_),
    .S(_01064_),
    .Y(_01099_)
  );
  OAI21X1 _07014_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01099_),
    .C(_01096_),
    .Y( execution_unit_0.alu_0.op_dst_6_ )
  );
  NAND2X1 _07015_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05690_),
    .Y(_01100_)
  );
  OAI21X1 _07016_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_7_ ),
    .Y(_01101_)
  );
  AOI22X1 _07017_ (
    .A(_01003_),
    .B(_01062_),
    .C(_01077_),
    .D(_01101_),
    .Y(_01102_)
  );
  MUX2X1 _07018_ (
    .A( execution_unit_0.inst_sext_7_ ),
    .B(_01102_),
    .S(_01064_),
    .Y(_01103_)
  );
  OAI21X1 _07019_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_01103_),
    .C(_01100_),
    .Y( execution_unit_0.alu_0.op_dst_7_ )
  );
  NAND2X1 _07020_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05691_),
    .Y(_01104_)
  );
  OAI21X1 _07021_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_8_ ),
    .Y(_01105_)
  );
  AOI22X1 _07022_ (
    .A(_00888_),
    .B(_01062_),
    .C(_01077_),
    .D(_01105_),
    .Y(_01106_)
  );
  NOR2X1 _07023_ (
    .A(_01064_),
    .B(_01106_),
    .Y(_01107_)
  );
  OAI21X1 _07024_ (
    .A( execution_unit_0.inst_sext_8_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01108_)
  );
  OAI21X1 _07025_ (
    .A(_01107_),
    .B(_01108_),
    .C(_01104_),
    .Y( execution_unit_0.alu_0.op_dst_8_ )
  );
  NAND2X1 _07026_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05692_),
    .Y(_01109_)
  );
  OAI21X1 _07027_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_9_ ),
    .Y(_01110_)
  );
  AOI22X1 _07028_ (
    .A(_00890_),
    .B(_01062_),
    .C(_01077_),
    .D(_01110_),
    .Y(_01111_)
  );
  NOR2X1 _07029_ (
    .A(_01064_),
    .B(_01111_),
    .Y(_01112_)
  );
  OAI21X1 _07030_ (
    .A( execution_unit_0.inst_sext_9_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01113_)
  );
  OAI21X1 _07031_ (
    .A(_01112_),
    .B(_01113_),
    .C(_01109_),
    .Y( execution_unit_0.alu_0.op_dst_9_ )
  );
  NAND2X1 _07032_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05678_),
    .Y(_01114_)
  );
  OAI21X1 _07033_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_10_ ),
    .Y(_01115_)
  );
  AOI22X1 _07034_ (
    .A(_00891_),
    .B(_01062_),
    .C(_01077_),
    .D(_01115_),
    .Y(_01116_)
  );
  NOR2X1 _07035_ (
    .A(_01064_),
    .B(_01116_),
    .Y(_01117_)
  );
  OAI21X1 _07036_ (
    .A( execution_unit_0.inst_sext_10_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01118_)
  );
  OAI21X1 _07037_ (
    .A(_01117_),
    .B(_01118_),
    .C(_01114_),
    .Y( execution_unit_0.alu_0.op_dst_10_ )
  );
  NAND2X1 _07038_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05679_),
    .Y(_01119_)
  );
  OAI21X1 _07039_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_11_ ),
    .Y(_01120_)
  );
  AOI22X1 _07040_ (
    .A(_00892_),
    .B(_01062_),
    .C(_01077_),
    .D(_01120_),
    .Y(_01121_)
  );
  NOR2X1 _07041_ (
    .A(_01064_),
    .B(_01121_),
    .Y(_01122_)
  );
  OAI21X1 _07042_ (
    .A( execution_unit_0.inst_sext_11_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01123_)
  );
  OAI21X1 _07043_ (
    .A(_01122_),
    .B(_01123_),
    .C(_01119_),
    .Y( execution_unit_0.alu_0.op_dst_11_ )
  );
  NAND2X1 _07044_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05680_),
    .Y(_01124_)
  );
  OAI21X1 _07045_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_12_ ),
    .Y(_01125_)
  );
  AOI22X1 _07046_ (
    .A(_00893_),
    .B(_01062_),
    .C(_01077_),
    .D(_01125_),
    .Y(_01126_)
  );
  NOR2X1 _07047_ (
    .A(_01064_),
    .B(_01126_),
    .Y(_01127_)
  );
  OAI21X1 _07048_ (
    .A( execution_unit_0.inst_sext_12_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01128_)
  );
  OAI21X1 _07049_ (
    .A(_01127_),
    .B(_01128_),
    .C(_01124_),
    .Y( execution_unit_0.alu_0.op_dst_12_ )
  );
  NAND2X1 _07050_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05681_),
    .Y(_01129_)
  );
  OAI21X1 _07051_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_13_ ),
    .Y(_01130_)
  );
  AOI22X1 _07052_ (
    .A(_00894_),
    .B(_01062_),
    .C(_01077_),
    .D(_01130_),
    .Y(_01131_)
  );
  NOR2X1 _07053_ (
    .A(_01064_),
    .B(_01131_),
    .Y(_01132_)
  );
  OAI21X1 _07054_ (
    .A( execution_unit_0.inst_sext_13_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01133_)
  );
  OAI21X1 _07055_ (
    .A(_01132_),
    .B(_01133_),
    .C(_01129_),
    .Y( execution_unit_0.alu_0.op_dst_13_ )
  );
  NAND2X1 _07056_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05682_),
    .Y(_01134_)
  );
  OAI21X1 _07057_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_14_ ),
    .Y(_01135_)
  );
  AOI22X1 _07058_ (
    .A(_00895_),
    .B(_01062_),
    .C(_01077_),
    .D(_01135_),
    .Y(_01136_)
  );
  NOR2X1 _07059_ (
    .A(_01064_),
    .B(_01136_),
    .Y(_01137_)
  );
  OAI21X1 _07060_ (
    .A( execution_unit_0.inst_sext_14_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01138_)
  );
  OAI21X1 _07061_ (
    .A(_01137_),
    .B(_01138_),
    .C(_01134_),
    .Y( execution_unit_0.alu_0.op_dst_14_ )
  );
  NAND2X1 _07062_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_05683_),
    .Y(_01139_)
  );
  OAI21X1 _07063_ (
    .A(_01053_),
    .B(_01056_),
    .C( dbg_0.dbg_reg_din_15_ ),
    .Y(_01140_)
  );
  AOI22X1 _07064_ (
    .A(_00896_),
    .B(_01062_),
    .C(_01077_),
    .D(_01140_),
    .Y(_01141_)
  );
  NOR2X1 _07065_ (
    .A(_01064_),
    .B(_01141_),
    .Y(_01142_)
  );
  OAI21X1 _07066_ (
    .A( execution_unit_0.inst_sext_15_ ),
    .B(_01065_),
    .C(_00905_),
    .Y(_01143_)
  );
  OAI21X1 _07067_ (
    .A(_01142_),
    .B(_01143_),
    .C(_01139_),
    .Y( execution_unit_0.alu_0.op_dst_15_ )
  );
  NAND2X1 _07068_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_0_ ),
    .Y(_01144_)
  );
  OAI21X1 _07069_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00906_),
    .C(_01144_),
    .Y( execution_unit_0.mdb_out_8_ )
  );
  NAND2X1 _07070_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_1_ ),
    .Y(_01145_)
  );
  OAI21X1 _07071_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00907_),
    .C(_01145_),
    .Y( execution_unit_0.mdb_out_9_ )
  );
  NAND2X1 _07072_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_2_ ),
    .Y(_01146_)
  );
  OAI21X1 _07073_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00908_),
    .C(_01146_),
    .Y( execution_unit_0.mdb_out_10_ )
  );
  NAND2X1 _07074_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_3_ ),
    .Y(_01147_)
  );
  OAI21X1 _07075_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00909_),
    .C(_01147_),
    .Y( execution_unit_0.mdb_out_11_ )
  );
  NAND2X1 _07076_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_4_ ),
    .Y(_01148_)
  );
  OAI21X1 _07077_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00910_),
    .C(_01148_),
    .Y( execution_unit_0.mdb_out_12_ )
  );
  NAND2X1 _07078_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_5_ ),
    .Y(_01149_)
  );
  OAI21X1 _07079_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00911_),
    .C(_01149_),
    .Y( execution_unit_0.mdb_out_13_ )
  );
  NAND2X1 _07080_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_6_ ),
    .Y(_01150_)
  );
  OAI21X1 _07081_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00912_),
    .C(_01150_),
    .Y( execution_unit_0.mdb_out_14_ )
  );
  NAND2X1 _07082_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( execution_unit_0.mdb_out_7_ ),
    .Y(_01151_)
  );
  OAI21X1 _07083_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00913_),
    .C(_01151_),
    .Y( execution_unit_0.mdb_out_15_ )
  );
  NAND3X1 _07084_ (
    .A( execution_unit_0.inst_as_0_ ),
    .B( execution_unit_0.inst_type_0_ ),
    .C(_01054_),
    .Y(_01152_)
  );
  NAND2X1 _07085_ (
    .A( execution_unit_0.inst_ad_0_ ),
    .B( execution_unit_0.inst_type_2_ ),
    .Y(_01153_)
  );
  OAI21X1 _07086_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_01153_),
    .C(_01152_),
    .Y(_01154_)
  );
  OAI21X1 _07087_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_01154_),
    .C( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01155_)
  );
  NAND2X1 _07088_ (
    .A(_00915_),
    .B(_01155_),
    .Y( execution_unit_0.reg_dest_wr )
  );
  NAND3X1 _07089_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_00916_),
    .C(_00921_),
    .Y(_01156_)
  );
  NAND2X1 _07090_ (
    .A(_00887_),
    .B(_01072_),
    .Y(_01157_)
  );
  OAI21X1 _07091_ (
    .A(_00933_),
    .B(_01157_),
    .C(_01156_),
    .Y(_01158_)
  );
  OR2X1 _07092_ (
    .A(_01074_),
    .B(_01158_),
    .Y( execution_unit_0.reg_sp_wr )
  );
  OAI21X1 _07093_ (
    .A(_00885_),
    .B(_00920_),
    .C(_01059_),
    .Y( execution_unit_0.reg_pc_call )
  );
  AOI22X1 _07094_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B( execution_unit_0.exec_done ),
    .C( execution_unit_0.alu_0.exec_cycle ),
    .D( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01159_)
  );
  OAI21X1 _07095_ (
    .A(_00886_),
    .B(_00926_),
    .C(_01159_),
    .Y( execution_unit_0.reg_incr )
  );
  AND2X1 _07096_ (
    .A(_00919_),
    .B(_00923_),
    .Y(_01160_)
  );
  OAI21X1 _07097_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_00942_),
    .C(_01156_),
    .Y(_01161_)
  );
  OAI21X1 _07098_ (
    .A(_01160_),
    .B(_01161_),
    .C(_00914_),
    .Y(_01162_)
  );
  OR2X1 _07099_ (
    .A( execution_unit_0.inst_type_0_ ),
    .B( execution_unit_0.inst_mov ),
    .Y(_01163_)
  );
  OAI22X1 _07100_ (
    .A(_00886_),
    .B(_00920_),
    .C(_00926_),
    .D( execution_unit_0.inst_as_5_ ),
    .Y(_01164_)
  );
  OAI21X1 _07101_ (
    .A(_00929_),
    .B(_01163_),
    .C(_01162_),
    .Y(_01165_)
  );
  OR2X1 _07102_ (
    .A(_01164_),
    .B(_01165_),
    .Y( dbg_0.UNUSED_eu_mb_en )
  );
  AOI21X1 _07103_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B( dbg_0.UNUSED_eu_mab_0_ ),
    .C(_01162_),
    .Y( dbg_0.UNUSED_eu_mb_wr_0_ )
  );
  AOI21X1 _07104_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_00917_),
    .C(_01162_),
    .Y( dbg_0.UNUSED_eu_mb_wr_1_ )
  );
  OAI21X1 _07105_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_00920_),
    .C(_00922_),
    .Y(_01166_)
  );
  NOR2X1 _07106_ (
    .A(_00928_),
    .B(_01166_),
    .Y(_01167_)
  );
  MUX2X1 _07107_ (
    .A( execution_unit_0.pc_nxt_0_ ),
    .B( execution_unit_0.alu_0.alu_out_0_ ),
    .S(_00928_),
    .Y(_01168_)
  );
  NAND2X1 _07108_ (
    .A( execution_unit_0.mdb_out_0_ ),
    .B(_01167_),
    .Y(_01169_)
  );
  OAI21X1 _07109_ (
    .A(_01167_),
    .B(_01168_),
    .C(_01169_),
    .Y(_00849_)
  );
  MUX2X1 _07110_ (
    .A( execution_unit_0.pc_nxt_1_ ),
    .B( execution_unit_0.alu_0.alu_out_1_ ),
    .S(_00928_),
    .Y(_01170_)
  );
  NAND2X1 _07111_ (
    .A( execution_unit_0.mdb_out_1_ ),
    .B(_01167_),
    .Y(_01171_)
  );
  OAI21X1 _07112_ (
    .A(_01167_),
    .B(_01170_),
    .C(_01171_),
    .Y(_00850_)
  );
  MUX2X1 _07113_ (
    .A( execution_unit_0.pc_nxt_2_ ),
    .B( execution_unit_0.alu_0.alu_out_2_ ),
    .S(_00928_),
    .Y(_01172_)
  );
  NAND2X1 _07114_ (
    .A( execution_unit_0.mdb_out_2_ ),
    .B(_01167_),
    .Y(_01173_)
  );
  OAI21X1 _07115_ (
    .A(_01167_),
    .B(_01172_),
    .C(_01173_),
    .Y(_00851_)
  );
  MUX2X1 _07116_ (
    .A( execution_unit_0.pc_nxt_3_ ),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .S(_00928_),
    .Y(_01174_)
  );
  NAND2X1 _07117_ (
    .A( execution_unit_0.mdb_out_3_ ),
    .B(_01167_),
    .Y(_01175_)
  );
  OAI21X1 _07118_ (
    .A(_01167_),
    .B(_01174_),
    .C(_01175_),
    .Y(_00852_)
  );
  MUX2X1 _07119_ (
    .A( execution_unit_0.pc_nxt_4_ ),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .S(_00928_),
    .Y(_01176_)
  );
  NAND2X1 _07120_ (
    .A( execution_unit_0.mdb_out_4_ ),
    .B(_01167_),
    .Y(_01177_)
  );
  OAI21X1 _07121_ (
    .A(_01167_),
    .B(_01176_),
    .C(_01177_),
    .Y(_00853_)
  );
  MUX2X1 _07122_ (
    .A( execution_unit_0.pc_nxt_5_ ),
    .B( execution_unit_0.alu_0.alu_out_5_ ),
    .S(_00928_),
    .Y(_01178_)
  );
  NAND2X1 _07123_ (
    .A( execution_unit_0.mdb_out_5_ ),
    .B(_01167_),
    .Y(_01179_)
  );
  OAI21X1 _07124_ (
    .A(_01167_),
    .B(_01178_),
    .C(_01179_),
    .Y(_00854_)
  );
  MUX2X1 _07125_ (
    .A( execution_unit_0.pc_nxt_6_ ),
    .B( execution_unit_0.alu_0.alu_out_6_ ),
    .S(_00928_),
    .Y(_01180_)
  );
  NAND2X1 _07126_ (
    .A( execution_unit_0.mdb_out_6_ ),
    .B(_01167_),
    .Y(_01181_)
  );
  OAI21X1 _07127_ (
    .A(_01167_),
    .B(_01180_),
    .C(_01181_),
    .Y(_00855_)
  );
  MUX2X1 _07128_ (
    .A( execution_unit_0.pc_nxt_7_ ),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .S(_00928_),
    .Y(_01182_)
  );
  NAND2X1 _07129_ (
    .A( execution_unit_0.mdb_out_7_ ),
    .B(_01167_),
    .Y(_01183_)
  );
  OAI21X1 _07130_ (
    .A(_01167_),
    .B(_01182_),
    .C(_01183_),
    .Y(_00856_)
  );
  MUX2X1 _07131_ (
    .A( execution_unit_0.pc_nxt_8_ ),
    .B( execution_unit_0.alu_0.alu_out_8_ ),
    .S(_00928_),
    .Y(_01184_)
  );
  NAND2X1 _07132_ (
    .A( execution_unit_0.mdb_out_nxt_8_ ),
    .B(_01167_),
    .Y(_01185_)
  );
  OAI21X1 _07133_ (
    .A(_01167_),
    .B(_01184_),
    .C(_01185_),
    .Y(_00857_)
  );
  MUX2X1 _07134_ (
    .A( execution_unit_0.pc_nxt_9_ ),
    .B( execution_unit_0.alu_0.alu_out_9_ ),
    .S(_00928_),
    .Y(_01186_)
  );
  NAND2X1 _07135_ (
    .A( execution_unit_0.mdb_out_nxt_9_ ),
    .B(_01167_),
    .Y(_01187_)
  );
  OAI21X1 _07136_ (
    .A(_01167_),
    .B(_01186_),
    .C(_01187_),
    .Y(_00858_)
  );
  MUX2X1 _07137_ (
    .A( execution_unit_0.pc_nxt_10_ ),
    .B( execution_unit_0.alu_0.alu_out_10_ ),
    .S(_00928_),
    .Y(_01188_)
  );
  NAND2X1 _07138_ (
    .A( execution_unit_0.mdb_out_nxt_10_ ),
    .B(_01167_),
    .Y(_01189_)
  );
  OAI21X1 _07139_ (
    .A(_01167_),
    .B(_01188_),
    .C(_01189_),
    .Y(_00859_)
  );
  MUX2X1 _07140_ (
    .A( execution_unit_0.pc_nxt_11_ ),
    .B( execution_unit_0.alu_0.alu_out_11_ ),
    .S(_00928_),
    .Y(_01190_)
  );
  NAND2X1 _07141_ (
    .A( execution_unit_0.mdb_out_nxt_11_ ),
    .B(_01167_),
    .Y(_01191_)
  );
  OAI21X1 _07142_ (
    .A(_01167_),
    .B(_01190_),
    .C(_01191_),
    .Y(_00860_)
  );
  MUX2X1 _07143_ (
    .A( execution_unit_0.pc_nxt_12_ ),
    .B( execution_unit_0.alu_0.alu_out_12_ ),
    .S(_00928_),
    .Y(_01192_)
  );
  NAND2X1 _07144_ (
    .A( execution_unit_0.mdb_out_nxt_12_ ),
    .B(_01167_),
    .Y(_01193_)
  );
  OAI21X1 _07145_ (
    .A(_01167_),
    .B(_01192_),
    .C(_01193_),
    .Y(_00861_)
  );
  MUX2X1 _07146_ (
    .A( execution_unit_0.pc_nxt_13_ ),
    .B( execution_unit_0.alu_0.alu_out_13_ ),
    .S(_00928_),
    .Y(_01194_)
  );
  NAND2X1 _07147_ (
    .A( execution_unit_0.mdb_out_nxt_13_ ),
    .B(_01167_),
    .Y(_01195_)
  );
  OAI21X1 _07148_ (
    .A(_01167_),
    .B(_01194_),
    .C(_01195_),
    .Y(_00862_)
  );
  MUX2X1 _07149_ (
    .A( execution_unit_0.pc_nxt_14_ ),
    .B( execution_unit_0.alu_0.alu_out_14_ ),
    .S(_00928_),
    .Y(_01196_)
  );
  NAND2X1 _07150_ (
    .A( execution_unit_0.mdb_out_nxt_14_ ),
    .B(_01167_),
    .Y(_01197_)
  );
  OAI21X1 _07151_ (
    .A(_01167_),
    .B(_01196_),
    .C(_01197_),
    .Y(_00863_)
  );
  MUX2X1 _07152_ (
    .A( execution_unit_0.pc_nxt_15_ ),
    .B( execution_unit_0.alu_0.alu_out_15_ ),
    .S(_00928_),
    .Y(_01198_)
  );
  NAND2X1 _07153_ (
    .A( execution_unit_0.mdb_out_nxt_15_ ),
    .B(_01167_),
    .Y(_01199_)
  );
  OAI21X1 _07154_ (
    .A(_01167_),
    .B(_01198_),
    .C(_01199_),
    .Y(_00864_)
  );
  NOR2X1 _07155_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_0_ ),
    .Y(_01200_)
  );
  AOI21X1 _07156_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00950_),
    .C(_01200_),
    .Y(_00865_)
  );
  NOR2X1 _07157_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_1_ ),
    .Y(_01201_)
  );
  AOI21X1 _07158_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00961_),
    .C(_01201_),
    .Y(_00866_)
  );
  NOR2X1 _07159_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_2_ ),
    .Y(_01202_)
  );
  AOI21X1 _07160_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00968_),
    .C(_01202_),
    .Y(_00867_)
  );
  NOR2X1 _07161_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_3_ ),
    .Y(_01203_)
  );
  AOI21X1 _07162_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00975_),
    .C(_01203_),
    .Y(_00868_)
  );
  NOR2X1 _07163_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_4_ ),
    .Y(_01204_)
  );
  AOI21X1 _07164_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00982_),
    .C(_01204_),
    .Y(_00869_)
  );
  NOR2X1 _07165_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_5_ ),
    .Y(_01205_)
  );
  AOI21X1 _07166_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00989_),
    .C(_01205_),
    .Y(_00870_)
  );
  NOR2X1 _07167_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_6_ ),
    .Y(_01206_)
  );
  AOI21X1 _07168_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00996_),
    .C(_01206_),
    .Y(_00871_)
  );
  NOR2X1 _07169_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_7_ ),
    .Y(_01207_)
  );
  AOI21X1 _07170_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_01003_),
    .C(_01207_),
    .Y(_00872_)
  );
  NAND2X1 _07171_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_8_ ),
    .Y(_01208_)
  );
  OAI21X1 _07172_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00897_),
    .C(_01208_),
    .Y(_00873_)
  );
  NAND2X1 _07173_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_9_ ),
    .Y(_01209_)
  );
  OAI21X1 _07174_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00898_),
    .C(_01209_),
    .Y(_00874_)
  );
  NAND2X1 _07175_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_10_ ),
    .Y(_01210_)
  );
  OAI21X1 _07176_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00899_),
    .C(_01210_),
    .Y(_00875_)
  );
  NAND2X1 _07177_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_11_ ),
    .Y(_01211_)
  );
  OAI21X1 _07178_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00900_),
    .C(_01211_),
    .Y(_00876_)
  );
  NAND2X1 _07179_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_12_ ),
    .Y(_01212_)
  );
  OAI21X1 _07180_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00901_),
    .C(_01212_),
    .Y(_00877_)
  );
  NAND2X1 _07181_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_13_ ),
    .Y(_01213_)
  );
  OAI21X1 _07182_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00902_),
    .C(_01213_),
    .Y(_00878_)
  );
  NAND2X1 _07183_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_14_ ),
    .Y(_01214_)
  );
  OAI21X1 _07184_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00903_),
    .C(_01214_),
    .Y(_00879_)
  );
  NAND2X1 _07185_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_15_ ),
    .Y(_01215_)
  );
  OAI21X1 _07186_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B(_00904_),
    .C(_01215_),
    .Y(_00880_)
  );
  OAI21X1 _07187_ (
    .A( execution_unit_0.mdb_in_buf_en ),
    .B( execution_unit_0.mdb_in_buf_valid ),
    .C(_00920_),
    .Y(_01216_)
  );
  INVX1 _07188_ (
    .A(_01216_),
    .Y(_00881_)
  );
  OAI21X1 _07189_ (
    .A(_01164_),
    .B(_01165_),
    .C( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01217_)
  );
  OAI21X1 _07190_ (
    .A(_00889_),
    .B( dbg_0.UNUSED_eu_mb_en ),
    .C(_01217_),
    .Y(_00882_)
  );
  DFFSR _07191_ (
    .CLK(dco_clk),
    .D(_00849_),
    .Q( execution_unit_0.mdb_out_0_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07192_ (
    .CLK(dco_clk),
    .D(_00850_),
    .Q( execution_unit_0.mdb_out_1_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07193_ (
    .CLK(dco_clk),
    .D(_00851_),
    .Q( execution_unit_0.mdb_out_2_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07194_ (
    .CLK(dco_clk),
    .D(_00852_),
    .Q( execution_unit_0.mdb_out_3_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07195_ (
    .CLK(dco_clk),
    .D(_00853_),
    .Q( execution_unit_0.mdb_out_4_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07196_ (
    .CLK(dco_clk),
    .D(_00854_),
    .Q( execution_unit_0.mdb_out_5_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07197_ (
    .CLK(dco_clk),
    .D(_00855_),
    .Q( execution_unit_0.mdb_out_6_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07198_ (
    .CLK(dco_clk),
    .D(_00856_),
    .Q( execution_unit_0.mdb_out_7_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07199_ (
    .CLK(dco_clk),
    .D(_00857_),
    .Q( execution_unit_0.mdb_out_nxt_8_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07200_ (
    .CLK(dco_clk),
    .D(_00858_),
    .Q( execution_unit_0.mdb_out_nxt_9_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07201_ (
    .CLK(dco_clk),
    .D(_00859_),
    .Q( execution_unit_0.mdb_out_nxt_10_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07202_ (
    .CLK(dco_clk),
    .D(_00860_),
    .Q( execution_unit_0.mdb_out_nxt_11_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07203_ (
    .CLK(dco_clk),
    .D(_00861_),
    .Q( execution_unit_0.mdb_out_nxt_12_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07204_ (
    .CLK(dco_clk),
    .D(_00862_),
    .Q( execution_unit_0.mdb_out_nxt_13_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07205_ (
    .CLK(dco_clk),
    .D(_00863_),
    .Q( execution_unit_0.mdb_out_nxt_14_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07206_ (
    .CLK(dco_clk),
    .D(_00864_),
    .Q( execution_unit_0.mdb_out_nxt_15_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07207_ (
    .CLK(dco_clk),
    .D(_00865_),
    .Q( execution_unit_0.mdb_in_buf_0_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07208_ (
    .CLK(dco_clk),
    .D(_00866_),
    .Q( execution_unit_0.mdb_in_buf_1_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07209_ (
    .CLK(dco_clk),
    .D(_00867_),
    .Q( execution_unit_0.mdb_in_buf_2_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07210_ (
    .CLK(dco_clk),
    .D(_00868_),
    .Q( execution_unit_0.mdb_in_buf_3_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07211_ (
    .CLK(dco_clk),
    .D(_00869_),
    .Q( execution_unit_0.mdb_in_buf_4_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07212_ (
    .CLK(dco_clk),
    .D(_00870_),
    .Q( execution_unit_0.mdb_in_buf_5_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07213_ (
    .CLK(dco_clk),
    .D(_00871_),
    .Q( execution_unit_0.mdb_in_buf_6_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07214_ (
    .CLK(dco_clk),
    .D(_00872_),
    .Q( execution_unit_0.mdb_in_buf_7_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07215_ (
    .CLK(dco_clk),
    .D(_00873_),
    .Q( execution_unit_0.mdb_in_buf_8_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07216_ (
    .CLK(dco_clk),
    .D(_00874_),
    .Q( execution_unit_0.mdb_in_buf_9_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07217_ (
    .CLK(dco_clk),
    .D(_00875_),
    .Q( execution_unit_0.mdb_in_buf_10_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07218_ (
    .CLK(dco_clk),
    .D(_00876_),
    .Q( execution_unit_0.mdb_in_buf_11_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07219_ (
    .CLK(dco_clk),
    .D(_00877_),
    .Q( execution_unit_0.mdb_in_buf_12_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07220_ (
    .CLK(dco_clk),
    .D(_00878_),
    .Q( execution_unit_0.mdb_in_buf_13_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07221_ (
    .CLK(dco_clk),
    .D(_00879_),
    .Q( execution_unit_0.mdb_in_buf_14_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07222_ (
    .CLK(dco_clk),
    .D(_00880_),
    .Q( execution_unit_0.mdb_in_buf_15_ ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07223_ (
    .CLK(dco_clk),
    .D(_00847_),
    .Q( execution_unit_0.mdb_in_buf_en ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07224_ (
    .CLK(dco_clk),
    .D(_00881_),
    .Q( execution_unit_0.mdb_in_buf_valid ),
    .R(_00848_),
    .S(1'h1)
  );
  DFFSR _07225_ (
    .CLK(dco_clk),
    .D(_00882_),
    .Q( execution_unit_0.mab_lsb ),
    .R(_00848_),
    .S(1'h1)
  );
  INVX1 _07226_ (
    .A( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01754_)
  );
  INVX1 _07227_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01218_)
  );
  INVX1 _07228_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01219_)
  );
  INVX1 _07229_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .Y(_01220_)
  );
  INVX1 _07230_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01221_)
  );
  INVX1 _07231_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .Y(_01222_)
  );
  INVX1 _07232_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01223_)
  );
  INVX1 _07233_ (
    .A( execution_unit_0.alu_0.inst_jmp_4_ ),
    .Y(_01224_)
  );
  INVX1 _07234_ (
    .A( execution_unit_0.alu_0.op_dst_3_ ),
    .Y(_01225_)
  );
  INVX1 _07235_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .Y(_01226_)
  );
  OR2X1 _07236_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B( execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_01227_)
  );
  NOR2X1 _07237_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01227_),
    .Y(_01228_)
  );
  OR2X1 _07238_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01227_),
    .Y(_01229_)
  );
  AOI21X1 _07239_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B( execution_unit_0.alu_0.inst_alu_2_ ),
    .C( execution_unit_0.alu_0.inst_alu_1_ ),
    .Y(_01230_)
  );
  NOR2X1 _07240_ (
    .A(_01754_),
    .B(_01230_),
    .Y(_01231_)
  );
  MUX2X1 _07241_ (
    .A( execution_unit_0.alu_0.inst_jmp_0_ ),
    .B( execution_unit_0.alu_0.inst_jmp_1_ ),
    .S( execution_unit_0.alu_0.status_1_ ),
    .Y(_01232_)
  );
  INVX1 _07242_ (
    .A(_01232_),
    .Y(_01233_)
  );
  MUX2X1 _07243_ (
    .A( execution_unit_0.alu_0.inst_jmp_2_ ),
    .B( execution_unit_0.alu_0.inst_jmp_3_ ),
    .S( execution_unit_0.alu_0.status_0_ ),
    .Y(_01234_)
  );
  OAI21X1 _07244_ (
    .A( execution_unit_0.alu_0.status_2_ ),
    .B(_01224_),
    .C(_01234_),
    .Y(_01235_)
  );
  NOR2X1 _07245_ (
    .A(_01233_),
    .B(_01235_),
    .Y(_01236_)
  );
  XOR2X1 _07246_ (
    .A( execution_unit_0.alu_0.status_3_ ),
    .B( execution_unit_0.alu_0.status_2_ ),
    .Y(_01237_)
  );
  MUX2X1 _07247_ (
    .A( execution_unit_0.alu_0.inst_jmp_5_ ),
    .B( execution_unit_0.alu_0.inst_jmp_6_ ),
    .S(_01237_),
    .Y(_01238_)
  );
  AND2X1 _07248_ (
    .A(_01236_),
    .B(_01238_),
    .Y(_01239_)
  );
  NAND2X1 _07249_ (
    .A(_01236_),
    .B(_01238_),
    .Y(_01240_)
  );
  NAND2X1 _07250_ (
    .A( execution_unit_0.alu_0.inst_alu_0_ ),
    .B( execution_unit_0.alu_0.exec_cycle ),
    .Y(_01241_)
  );
  XNOR2X1 _07251_ (
    .A( execution_unit_0.alu_0.alu_swpb_8_ ),
    .B(_01241_),
    .Y(_01242_)
  );
  NOR2X1 _07252_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01242_),
    .Y(_01243_)
  );
  OR2X1 _07253_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01242_),
    .Y(_01244_)
  );
  AND2X1 _07254_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01242_),
    .Y(_01245_)
  );
  NAND2X1 _07255_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01242_),
    .Y(_01246_)
  );
  NAND2X1 _07256_ (
    .A(_01239_),
    .B(_01246_),
    .Y(_01247_)
  );
  OAI21X1 _07257_ (
    .A( execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01239_),
    .C(_01244_),
    .Y(_01248_)
  );
  AOI21X1 _07258_ (
    .A(_01239_),
    .B(_01245_),
    .C(_01248_),
    .Y( dbg_0.UNUSED_eu_mab_0_ )
  );
  NAND2X1 _07259_ (
    .A(_01231_),
    .B( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01249_)
  );
  XNOR2X1 _07260_ (
    .A(_01231_),
    .B( dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01250_)
  );
  NAND2X1 _07261_ (
    .A(_01244_),
    .B(_01246_),
    .Y(_01251_)
  );
  OR2X1 _07262_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.inst_so_3_ ),
    .Y(_01252_)
  );
  NOR2X1 _07263_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01253_)
  );
  NAND3X1 _07264_ (
    .A(_01220_),
    .B(_01221_),
    .C(_01253_),
    .Y(_01254_)
  );
  NOR2X1 _07265_ (
    .A(_01252_),
    .B(_01254_),
    .Y(_01255_)
  );
  AOI21X1 _07266_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_swpb_0_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01256_)
  );
  AOI22X1 _07267_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B( execution_unit_0.alu_0.inst_alu_10_ ),
    .C( execution_unit_0.alu_0.inst_so_3_ ),
    .D( execution_unit_0.alu_0.alu_swpb_8_ ),
    .Y(_01257_)
  );
  NAND2X1 _07268_ (
    .A(_01256_),
    .B(_01257_),
    .Y(_01258_)
  );
  AOI21X1 _07269_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01244_),
    .C(_01258_),
    .Y(_01259_)
  );
  AOI22X1 _07270_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01245_),
    .C(_01255_),
    .D(_01242_),
    .Y(_01260_)
  );
  AND2X1 _07271_ (
    .A(_01259_),
    .B(_01260_),
    .Y(_01261_)
  );
  OAI21X1 _07272_ (
    .A(_01220_),
    .B(_01251_),
    .C(_01261_),
    .Y(_01262_)
  );
  XNOR2X1 _07273_ (
    .A(_01222_),
    .B(_01251_),
    .Y(_01263_)
  );
  AOI21X1 _07274_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01263_),
    .C(_01229_),
    .Y(_01264_)
  );
  NAND2X1 _07275_ (
    .A(_01262_),
    .B(_01264_),
    .Y(_01265_)
  );
  OAI21X1 _07276_ (
    .A(_01228_),
    .B(_01250_),
    .C(_01265_),
    .Y( execution_unit_0.alu_0.alu_out_0_ )
  );
  XNOR2X1 _07277_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B(_01241_),
    .Y(_01266_)
  );
  NOR2X1 _07278_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01266_),
    .Y(_01267_)
  );
  AND2X1 _07279_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01266_),
    .Y(_01268_)
  );
  INVX1 _07280_ (
    .A(_01268_),
    .Y(_01269_)
  );
  NOR2X1 _07281_ (
    .A(_01267_),
    .B(_01268_),
    .Y(_01270_)
  );
  XNOR2X1 _07282_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01266_),
    .Y(_01271_)
  );
  NAND2X1 _07283_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01240_),
    .Y(_01272_)
  );
  NOR2X1 _07284_ (
    .A(_01246_),
    .B(_01271_),
    .Y(_01273_)
  );
  OAI21X1 _07285_ (
    .A(_01240_),
    .B(_01273_),
    .C(_01272_),
    .Y(_01274_)
  );
  OAI21X1 _07286_ (
    .A(_01247_),
    .B(_01270_),
    .C(_01274_),
    .Y(_01275_)
  );
  INVX1 _07287_ (
    .A(_01275_),
    .Y( dbg_0.UNUSED_eu_mab_1_ )
  );
  NOR2X1 _07288_ (
    .A(_01249_),
    .B(_01275_),
    .Y(_01276_)
  );
  NAND2X1 _07289_ (
    .A(_01249_),
    .B(_01275_),
    .Y(_01277_)
  );
  OAI21X1 _07290_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01227_),
    .C(_01277_),
    .Y(_01278_)
  );
  AOI21X1 _07291_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B(_01244_),
    .C(_01245_),
    .Y(_01279_)
  );
  OAI21X1 _07292_ (
    .A(_01222_),
    .B(_01243_),
    .C(_01246_),
    .Y(_01280_)
  );
  XNOR2X1 _07293_ (
    .A(_01270_),
    .B(_01279_),
    .Y(_01281_)
  );
  INVX1 _07294_ (
    .A(_01281_),
    .Y(_01282_)
  );
  XNOR2X1 _07295_ (
    .A( execution_unit_0.alu_0.alu_shift_2_ ),
    .B(_01241_),
    .Y(_01283_)
  );
  INVX1 _07296_ (
    .A(_01283_),
    .Y(_01284_)
  );
  NAND2X1 _07297_ (
    .A( execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01283_),
    .Y(_01285_)
  );
  INVX1 _07298_ (
    .A(_01285_),
    .Y(_01286_)
  );
  NAND2X1 _07299_ (
    .A(_01225_),
    .B(_01284_),
    .Y(_01287_)
  );
  NAND2X1 _07300_ (
    .A(_01285_),
    .B(_01287_),
    .Y(_01288_)
  );
  XNOR2X1 _07301_ (
    .A( execution_unit_0.alu_0.alu_shift_1_ ),
    .B(_01241_),
    .Y(_01289_)
  );
  AND2X1 _07302_ (
    .A( execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01289_),
    .Y(_01290_)
  );
  INVX1 _07303_ (
    .A(_01290_),
    .Y(_01291_)
  );
  AOI21X1 _07304_ (
    .A(_01270_),
    .B(_01280_),
    .C(_01268_),
    .Y(_01292_)
  );
  OAI21X1 _07305_ (
    .A(_01271_),
    .B(_01279_),
    .C(_01269_),
    .Y(_01293_)
  );
  NOR2X1 _07306_ (
    .A( execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01289_),
    .Y(_01294_)
  );
  INVX1 _07307_ (
    .A(_01294_),
    .Y(_01295_)
  );
  NAND2X1 _07308_ (
    .A(_01291_),
    .B(_01295_),
    .Y(_01296_)
  );
  AOI21X1 _07309_ (
    .A(_01293_),
    .B(_01295_),
    .C(_01290_),
    .Y(_01297_)
  );
  OAI21X1 _07310_ (
    .A(_01292_),
    .B(_01294_),
    .C(_01291_),
    .Y(_01298_)
  );
  AOI21X1 _07311_ (
    .A(_01287_),
    .B(_01298_),
    .C(_01286_),
    .Y(_01299_)
  );
  OAI21X1 _07312_ (
    .A(_01288_),
    .B(_01297_),
    .C(_01285_),
    .Y(_01300_)
  );
  XNOR2X1 _07313_ (
    .A(_01288_),
    .B(_01298_),
    .Y(_01301_)
  );
  XNOR2X1 _07314_ (
    .A(_01288_),
    .B(_01297_),
    .Y(_01302_)
  );
  XNOR2X1 _07315_ (
    .A(_01292_),
    .B(_01296_),
    .Y(_01303_)
  );
  AND2X1 _07316_ (
    .A(_01282_),
    .B(_01303_),
    .Y(_01304_)
  );
  NAND2X1 _07317_ (
    .A(_01282_),
    .B(_01303_),
    .Y(_01305_)
  );
  AOI21X1 _07318_ (
    .A(_01301_),
    .B(_01305_),
    .C(_01300_),
    .Y(_01306_)
  );
  OAI21X1 _07319_ (
    .A(_01302_),
    .B(_01304_),
    .C(_01299_),
    .Y(_01307_)
  );
  NOR2X1 _07320_ (
    .A(_01281_),
    .B(_01306_),
    .Y(_01308_)
  );
  OAI21X1 _07321_ (
    .A(_01282_),
    .B(_01307_),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01309_)
  );
  OAI21X1 _07322_ (
    .A( execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01266_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01310_)
  );
  AOI22X1 _07323_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B( execution_unit_0.alu_0.inst_so_3_ ),
    .C( execution_unit_0.alu_0.alu_shift_1_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01311_)
  );
  NAND2X1 _07324_ (
    .A(_01223_),
    .B(_01311_),
    .Y(_01312_)
  );
  AOI21X1 _07325_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_8_ ),
    .C(_01312_),
    .Y(_01313_)
  );
  AOI22X1 _07326_ (
    .A(_01255_),
    .B(_01266_),
    .C(_01268_),
    .D( execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01314_)
  );
  NAND3X1 _07327_ (
    .A(_01310_),
    .B(_01313_),
    .C(_01314_),
    .Y(_01315_)
  );
  AOI21X1 _07328_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01270_),
    .C(_01315_),
    .Y(_01316_)
  );
  NOR2X1 _07329_ (
    .A(_01229_),
    .B(_01316_),
    .Y(_01317_)
  );
  OAI21X1 _07330_ (
    .A(_01308_),
    .B(_01309_),
    .C(_01317_),
    .Y(_01318_)
  );
  OAI21X1 _07331_ (
    .A(_01276_),
    .B(_01278_),
    .C(_01318_),
    .Y( execution_unit_0.alu_0.alu_out_1_ )
  );
  AOI21X1 _07332_ (
    .A(_01239_),
    .B(_01290_),
    .C(_01294_),
    .Y(_01319_)
  );
  OAI21X1 _07333_ (
    .A( execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01239_),
    .C(_01319_),
    .Y(_01320_)
  );
  OAI21X1 _07334_ (
    .A(_01268_),
    .B(_01273_),
    .C(_01239_),
    .Y(_01321_)
  );
  XOR2X1 _07335_ (
    .A(_01320_),
    .B(_01321_),
    .Y( dbg_0.UNUSED_eu_mab_2_ )
  );
  NAND2X1 _07336_ (
    .A(_01276_),
    .B( dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_01322_)
  );
  XNOR2X1 _07337_ (
    .A(_01276_),
    .B( dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_01323_)
  );
  NAND2X1 _07338_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01228_),
    .Y(_01324_)
  );
  NAND2X1 _07339_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_1_ ),
    .Y(_01325_)
  );
  AOI22X1 _07340_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_2_ ),
    .C( execution_unit_0.alu_0.alu_shift_9_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01326_)
  );
  NAND3X1 _07341_ (
    .A(_01228_),
    .B(_01325_),
    .C(_01326_),
    .Y(_01327_)
  );
  AOI21X1 _07342_ (
    .A(_01255_),
    .B(_01289_),
    .C(_01327_),
    .Y(_01328_)
  );
  OAI21X1 _07343_ (
    .A(_01219_),
    .B(_01294_),
    .C(_01328_),
    .Y(_01329_)
  );
  AOI21X1 _07344_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01290_),
    .C(_01329_),
    .Y(_01330_)
  );
  OAI21X1 _07345_ (
    .A(_01220_),
    .B(_01296_),
    .C(_01330_),
    .Y(_01331_)
  );
  XNOR2X1 _07346_ (
    .A(_01303_),
    .B(_01308_),
    .Y(_01332_)
  );
  AOI22X1 _07347_ (
    .A(_01324_),
    .B(_01331_),
    .C(_01332_),
    .D( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01333_)
  );
  AOI21X1 _07348_ (
    .A(_01229_),
    .B(_01323_),
    .C(_01333_),
    .Y( execution_unit_0.alu_0.alu_out_2_ )
  );
  OAI22X1 _07349_ (
    .A(_01240_),
    .B(_01291_),
    .C(_01296_),
    .D(_01321_),
    .Y(_01334_)
  );
  OAI21X1 _07350_ (
    .A(_01240_),
    .B(_01284_),
    .C(_01225_),
    .Y(_01335_)
  );
  OAI21X1 _07351_ (
    .A(_01240_),
    .B(_01285_),
    .C(_01335_),
    .Y(_01336_)
  );
  XOR2X1 _07352_ (
    .A(_01334_),
    .B(_01336_),
    .Y(_01337_)
  );
  INVX1 _07353_ (
    .A(_01337_),
    .Y( dbg_0.UNUSED_eu_mab_3_ )
  );
  NOR2X1 _07354_ (
    .A(_01322_),
    .B(_01337_),
    .Y(_01338_)
  );
  XNOR2X1 _07355_ (
    .A(_01322_),
    .B(_01337_),
    .Y(_01339_)
  );
  OAI21X1 _07356_ (
    .A(_01299_),
    .B(_01304_),
    .C(_01302_),
    .Y(_01340_)
  );
  AND2X1 _07357_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01340_),
    .Y(_01341_)
  );
  OAI21X1 _07358_ (
    .A(_01302_),
    .B(_01304_),
    .C(_01341_),
    .Y(_01342_)
  );
  OAI21X1 _07359_ (
    .A( execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01283_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01343_)
  );
  AOI22X1 _07360_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_2_ ),
    .C( execution_unit_0.alu_0.alu_shift_3_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01344_)
  );
  AOI22X1 _07361_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_10_ ),
    .C(_01255_),
    .D(_01283_),
    .Y(_01345_)
  );
  OAI21X1 _07362_ (
    .A(_01218_),
    .B(_01285_),
    .C(_01345_),
    .Y(_01346_)
  );
  INVX1 _07363_ (
    .A(_01346_),
    .Y(_01347_)
  );
  NAND3X1 _07364_ (
    .A(_01343_),
    .B(_01344_),
    .C(_01347_),
    .Y(_01348_)
  );
  OAI21X1 _07365_ (
    .A(_01220_),
    .B(_01288_),
    .C(_01228_),
    .Y(_01349_)
  );
  OAI21X1 _07366_ (
    .A(_01348_),
    .B(_01349_),
    .C(_01324_),
    .Y(_01350_)
  );
  AOI22X1 _07367_ (
    .A(_01229_),
    .B(_01339_),
    .C(_01342_),
    .D(_01350_),
    .Y( execution_unit_0.alu_0.alu_out_3_ )
  );
  XNOR2X1 _07368_ (
    .A( execution_unit_0.alu_0.alu_shift_3_ ),
    .B(_01241_),
    .Y(_01351_)
  );
  AND2X1 _07369_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01351_),
    .Y(_01352_)
  );
  NAND2X1 _07370_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01351_),
    .Y(_01353_)
  );
  NAND2X1 _07371_ (
    .A(_01239_),
    .B(_01351_),
    .Y(_01354_)
  );
  XOR2X1 _07372_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01354_),
    .Y(_01355_)
  );
  AOI22X1 _07373_ (
    .A(_01239_),
    .B(_01286_),
    .C(_01334_),
    .D(_01335_),
    .Y(_01356_)
  );
  XOR2X1 _07374_ (
    .A(_01355_),
    .B(_01356_),
    .Y( dbg_0.UNUSED_eu_mab_4_ )
  );
  NOR2X1 _07375_ (
    .A( execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01351_),
    .Y(_01357_)
  );
  NOR2X1 _07376_ (
    .A(_01352_),
    .B(_01357_),
    .Y(_01358_)
  );
  INVX1 _07377_ (
    .A(_01358_),
    .Y(_01359_)
  );
  NOR3X1 _07378_ (
    .A(_01299_),
    .B(_01302_),
    .C(_01304_),
    .Y(_01360_)
  );
  NAND3X1 _07379_ (
    .A(_01300_),
    .B(_01301_),
    .C(_01305_),
    .Y(_01361_)
  );
  OAI21X1 _07380_ (
    .A(_01306_),
    .B(_01360_),
    .C(_01359_),
    .Y(_01362_)
  );
  NOR3X1 _07381_ (
    .A(_01306_),
    .B(_01359_),
    .C(_01360_),
    .Y(_01363_)
  );
  NAND3X1 _07382_ (
    .A(_01307_),
    .B(_01358_),
    .C(_01361_),
    .Y(_01364_)
  );
  AND2X1 _07383_ (
    .A(_01362_),
    .B(_01364_),
    .Y(_01365_)
  );
  NAND2X1 _07384_ (
    .A(_01338_),
    .B( dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_01366_)
  );
  XNOR2X1 _07385_ (
    .A(_01338_),
    .B( dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_01367_)
  );
  AOI21X1 _07386_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_3_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01368_)
  );
  AOI22X1 _07387_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_4_ ),
    .C( execution_unit_0.alu_0.alu_shift_11_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01369_)
  );
  NAND3X1 _07388_ (
    .A(_01228_),
    .B(_01368_),
    .C(_01369_),
    .Y(_01370_)
  );
  AOI21X1 _07389_ (
    .A(_01255_),
    .B(_01351_),
    .C(_01370_),
    .Y(_01371_)
  );
  OAI21X1 _07390_ (
    .A(_01219_),
    .B(_01357_),
    .C(_01371_),
    .Y(_01372_)
  );
  AOI21X1 _07391_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01352_),
    .C(_01372_),
    .Y(_01373_)
  );
  OAI21X1 _07392_ (
    .A(_01220_),
    .B(_01359_),
    .C(_01373_),
    .Y(_01374_)
  );
  OAI21X1 _07393_ (
    .A(_01324_),
    .B(_01365_),
    .C(_01374_),
    .Y(_01375_)
  );
  AOI21X1 _07394_ (
    .A(_01229_),
    .B(_01367_),
    .C(_01375_),
    .Y( execution_unit_0.alu_0.alu_out_4_ )
  );
  OAI22X1 _07395_ (
    .A(_01240_),
    .B(_01353_),
    .C(_01355_),
    .D(_01356_),
    .Y(_01376_)
  );
  INVX1 _07396_ (
    .A(_01376_),
    .Y(_01377_)
  );
  XNOR2X1 _07397_ (
    .A( execution_unit_0.alu_0.alu_shift_4_ ),
    .B(_01241_),
    .Y(_01378_)
  );
  AND2X1 _07398_ (
    .A( execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01378_),
    .Y(_01379_)
  );
  NAND2X1 _07399_ (
    .A( execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01378_),
    .Y(_01380_)
  );
  NOR2X1 _07400_ (
    .A(_01240_),
    .B(_01380_),
    .Y(_01381_)
  );
  AOI21X1 _07401_ (
    .A(_01239_),
    .B(_01378_),
    .C( execution_unit_0.alu_0.op_dst_5_ ),
    .Y(_01382_)
  );
  OR2X1 _07402_ (
    .A(_01381_),
    .B(_01382_),
    .Y(_01383_)
  );
  NOR2X1 _07403_ (
    .A(_01377_),
    .B(_01383_),
    .Y(_01384_)
  );
  XOR2X1 _07404_ (
    .A(_01376_),
    .B(_01383_),
    .Y(_01385_)
  );
  INVX1 _07405_ (
    .A(_01385_),
    .Y( dbg_0.UNUSED_eu_mab_5_ )
  );
  NOR2X1 _07406_ (
    .A(_01366_),
    .B(_01385_),
    .Y(_01386_)
  );
  INVX1 _07407_ (
    .A(_01386_),
    .Y(_01387_)
  );
  AOI21X1 _07408_ (
    .A(_01366_),
    .B(_01385_),
    .C(_01228_),
    .Y(_01388_)
  );
  OR2X1 _07409_ (
    .A( execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01378_),
    .Y(_01389_)
  );
  AND2X1 _07410_ (
    .A(_01380_),
    .B(_01389_),
    .Y(_01390_)
  );
  NAND2X1 _07411_ (
    .A(_01380_),
    .B(_01389_),
    .Y(_01391_)
  );
  AOI21X1 _07412_ (
    .A(_01353_),
    .B(_01364_),
    .C(_01391_),
    .Y(_01392_)
  );
  OAI21X1 _07413_ (
    .A(_01352_),
    .B(_01363_),
    .C(_01390_),
    .Y(_01393_)
  );
  NAND3X1 _07414_ (
    .A(_01353_),
    .B(_01364_),
    .C(_01391_),
    .Y(_01394_)
  );
  NAND2X1 _07415_ (
    .A(_01393_),
    .B(_01394_),
    .Y(_01395_)
  );
  XNOR2X1 _07416_ (
    .A( execution_unit_0.alu_0.alu_shift_5_ ),
    .B(_01241_),
    .Y(_01396_)
  );
  AND2X1 _07417_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01396_),
    .Y(_01397_)
  );
  NAND2X1 _07418_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01396_),
    .Y(_01398_)
  );
  XNOR2X1 _07419_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01396_),
    .Y(_01399_)
  );
  INVX1 _07420_ (
    .A(_01399_),
    .Y(_01400_)
  );
  NOR2X1 _07421_ (
    .A(_01379_),
    .B(_01392_),
    .Y(_01401_)
  );
  AOI21X1 _07422_ (
    .A(_01380_),
    .B(_01393_),
    .C(_01399_),
    .Y(_01402_)
  );
  OAI21X1 _07423_ (
    .A(_01379_),
    .B(_01392_),
    .C(_01400_),
    .Y(_01403_)
  );
  XNOR2X1 _07424_ (
    .A(_01399_),
    .B(_01401_),
    .Y(_01404_)
  );
  NAND2X1 _07425_ (
    .A(_01395_),
    .B(_01404_),
    .Y(_01405_)
  );
  OAI21X1 _07426_ (
    .A(_01399_),
    .B(_01401_),
    .C(_01398_),
    .Y(_01406_)
  );
  XNOR2X1 _07427_ (
    .A( execution_unit_0.alu_0.alu_shift_6_ ),
    .B(_01241_),
    .Y(_01407_)
  );
  AND2X1 _07428_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01407_),
    .Y(_01408_)
  );
  NAND2X1 _07429_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01407_),
    .Y(_01409_)
  );
  OR2X1 _07430_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01407_),
    .Y(_01410_)
  );
  NAND2X1 _07431_ (
    .A(_01409_),
    .B(_01410_),
    .Y(_01411_)
  );
  INVX1 _07432_ (
    .A(_01411_),
    .Y(_01412_)
  );
  NAND3X1 _07433_ (
    .A(_01398_),
    .B(_01403_),
    .C(_01412_),
    .Y(_01413_)
  );
  OAI21X1 _07434_ (
    .A(_01397_),
    .B(_01402_),
    .C(_01411_),
    .Y(_01414_)
  );
  NAND2X1 _07435_ (
    .A(_01413_),
    .B(_01414_),
    .Y(_01415_)
  );
  AOI22X1 _07436_ (
    .A(_01395_),
    .B(_01404_),
    .C(_01413_),
    .D(_01414_),
    .Y(_01416_)
  );
  NAND2X1 _07437_ (
    .A(_01405_),
    .B(_01415_),
    .Y(_01417_)
  );
  OAI21X1 _07438_ (
    .A(_01406_),
    .B(_01408_),
    .C(_01410_),
    .Y(_01418_)
  );
  NAND2X1 _07439_ (
    .A(_01417_),
    .B(_01418_),
    .Y(_01419_)
  );
  NAND2X1 _07440_ (
    .A(_01395_),
    .B(_01419_),
    .Y(_01420_)
  );
  XOR2X1 _07441_ (
    .A(_01395_),
    .B(_01419_),
    .Y(_01421_)
  );
  AOI21X1 _07442_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_5_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01422_)
  );
  AOI22X1 _07443_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_4_ ),
    .C( execution_unit_0.alu_0.alu_shift_12_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01423_)
  );
  NAND2X1 _07444_ (
    .A(_01422_),
    .B(_01423_),
    .Y(_01424_)
  );
  AOI21X1 _07445_ (
    .A(_01255_),
    .B(_01378_),
    .C(_01424_),
    .Y(_01425_)
  );
  OAI21X1 _07446_ (
    .A(_01218_),
    .B(_01380_),
    .C(_01425_),
    .Y(_01426_)
  );
  AOI21X1 _07447_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01389_),
    .C(_01426_),
    .Y(_01427_)
  );
  OAI21X1 _07448_ (
    .A(_01220_),
    .B(_01391_),
    .C(_01427_),
    .Y(_01428_)
  );
  NAND2X1 _07449_ (
    .A(_01228_),
    .B(_01428_),
    .Y(_01429_)
  );
  AOI21X1 _07450_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01421_),
    .C(_01429_),
    .Y(_01430_)
  );
  AOI21X1 _07451_ (
    .A(_01387_),
    .B(_01388_),
    .C(_01430_),
    .Y(_01431_)
  );
  INVX1 _07452_ (
    .A(_01431_),
    .Y( execution_unit_0.alu_0.alu_out_5_ )
  );
  NOR2X1 _07453_ (
    .A(_01381_),
    .B(_01384_),
    .Y(_01432_)
  );
  NOR2X1 _07454_ (
    .A(_01240_),
    .B(_01398_),
    .Y(_01433_)
  );
  AOI21X1 _07455_ (
    .A(_01239_),
    .B(_01396_),
    .C( execution_unit_0.alu_0.op_dst_6_ ),
    .Y(_01434_)
  );
  OR2X1 _07456_ (
    .A(_01433_),
    .B(_01434_),
    .Y(_01435_)
  );
  OAI21X1 _07457_ (
    .A(_01433_),
    .B(_01434_),
    .C(_01432_),
    .Y(_01436_)
  );
  OR2X1 _07458_ (
    .A(_01432_),
    .B(_01435_),
    .Y(_01437_)
  );
  NAND2X1 _07459_ (
    .A(_01436_),
    .B(_01437_),
    .Y(_01438_)
  );
  INVX1 _07460_ (
    .A(_01438_),
    .Y( dbg_0.UNUSED_eu_mab_6_ )
  );
  NOR2X1 _07461_ (
    .A(_01387_),
    .B(_01438_),
    .Y(_01439_)
  );
  XOR2X1 _07462_ (
    .A(_01386_),
    .B(_01438_),
    .Y(_01440_)
  );
  OAI21X1 _07463_ (
    .A( execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01396_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01441_)
  );
  NAND2X1 _07464_ (
    .A(_01255_),
    .B(_01396_),
    .Y(_01442_)
  );
  AOI22X1 _07465_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_5_ ),
    .C( execution_unit_0.alu_0.alu_shift_13_ ),
    .D( execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01443_)
  );
  NAND2X1 _07466_ (
    .A(_01228_),
    .B(_01443_),
    .Y(_01444_)
  );
  AOI21X1 _07467_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_6_ ),
    .C(_01444_),
    .Y(_01445_)
  );
  NAND2X1 _07468_ (
    .A(_01441_),
    .B(_01442_),
    .Y(_01446_)
  );
  OAI21X1 _07469_ (
    .A(_01220_),
    .B(_01399_),
    .C(_01445_),
    .Y(_01447_)
  );
  NOR2X1 _07470_ (
    .A(_01446_),
    .B(_01447_),
    .Y(_01448_)
  );
  OAI21X1 _07471_ (
    .A(_01218_),
    .B(_01398_),
    .C(_01448_),
    .Y(_01449_)
  );
  XOR2X1 _07472_ (
    .A(_01404_),
    .B(_01420_),
    .Y(_01450_)
  );
  AOI22X1 _07473_ (
    .A(_01324_),
    .B(_01449_),
    .C(_01450_),
    .D( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01451_)
  );
  AOI21X1 _07474_ (
    .A(_01229_),
    .B(_01440_),
    .C(_01451_),
    .Y( execution_unit_0.alu_0.alu_out_6_ )
  );
  AOI21X1 _07475_ (
    .A(_01405_),
    .B(_01410_),
    .C(_01415_),
    .Y(_01452_)
  );
  NOR2X1 _07476_ (
    .A(_01416_),
    .B(_01452_),
    .Y(_01453_)
  );
  OAI21X1 _07477_ (
    .A(_01240_),
    .B(_01398_),
    .C(_01437_),
    .Y(_01454_)
  );
  NOR2X1 _07478_ (
    .A(_01240_),
    .B(_01409_),
    .Y(_01455_)
  );
  OAI21X1 _07479_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01239_),
    .C(_01410_),
    .Y(_01456_)
  );
  NOR2X1 _07480_ (
    .A(_01455_),
    .B(_01456_),
    .Y(_01457_)
  );
  XOR2X1 _07481_ (
    .A(_01454_),
    .B(_01457_),
    .Y( dbg_0.UNUSED_eu_mab_7_ )
  );
  NAND2X1 _07482_ (
    .A(_01439_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01458_)
  );
  XNOR2X1 _07483_ (
    .A(_01439_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01459_)
  );
  OAI21X1 _07484_ (
    .A(_01220_),
    .B(_01408_),
    .C(_01219_),
    .Y(_01460_)
  );
  OAI21X1 _07485_ (
    .A( execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01407_),
    .C(_01460_),
    .Y(_01461_)
  );
  MUX2X1 _07486_ (
    .A( execution_unit_0.alu_0.alu_shift_6_ ),
    .B( execution_unit_0.alu_0.alu_shift_14_ ),
    .S( execution_unit_0.alu_0.inst_bw ),
    .Y(_01462_)
  );
  NOR2X1 _07487_ (
    .A( execution_unit_0.alu_0.inst_so_0_ ),
    .B(_01462_),
    .Y(_01463_)
  );
  AOI21X1 _07488_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B( execution_unit_0.alu_0.inst_so_0_ ),
    .C(_01463_),
    .Y(_01464_)
  );
  OAI21X1 _07489_ (
    .A( execution_unit_0.alu_0.alu_swpb_0_ ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .C( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01465_)
  );
  AOI21X1 _07490_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_01464_),
    .C(_01465_),
    .Y(_01466_)
  );
  AOI21X1 _07491_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_6_ ),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01467_)
  );
  AOI21X1 _07492_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_14_ ),
    .C(_01229_),
    .Y(_01468_)
  );
  NAND2X1 _07493_ (
    .A(_01467_),
    .B(_01468_),
    .Y(_01469_)
  );
  AOI21X1 _07494_ (
    .A(_01255_),
    .B(_01407_),
    .C(_01469_),
    .Y(_01470_)
  );
  OAI21X1 _07495_ (
    .A(_01218_),
    .B(_01409_),
    .C(_01470_),
    .Y(_01471_)
  );
  NOR2X1 _07496_ (
    .A(_01466_),
    .B(_01471_),
    .Y(_01472_)
  );
  AOI22X1 _07497_ (
    .A(_01229_),
    .B(_01459_),
    .C(_01461_),
    .D(_01472_),
    .Y(_01473_)
  );
  OAI21X1 _07498_ (
    .A(_01324_),
    .B(_01453_),
    .C(_01473_),
    .Y(_01474_)
  );
  INVX1 _07499_ (
    .A(_01474_),
    .Y( execution_unit_0.alu_0.alu_out_7_ )
  );
  AOI21X1 _07500_ (
    .A(_01410_),
    .B(_01433_),
    .C(_01455_),
    .Y(_01475_)
  );
  OAI21X1 _07501_ (
    .A(_01437_),
    .B(_01456_),
    .C(_01475_),
    .Y(_01476_)
  );
  NOR2X1 _07502_ (
    .A(_01754_),
    .B(_01226_),
    .Y(_01477_)
  );
  NAND2X1 _07503_ (
    .A( execution_unit_0.alu_0.exec_cycle ),
    .B( execution_unit_0.alu_0.inst_bw ),
    .Y(_01478_)
  );
  XOR2X1 _07504_ (
    .A( execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(_01241_),
    .Y(_01479_)
  );
  NOR2X1 _07505_ (
    .A(_01477_),
    .B(_01479_),
    .Y(_01480_)
  );
  OAI21X1 _07506_ (
    .A(_01754_),
    .B(_01226_),
    .C( execution_unit_0.alu_0.op_dst_8_ ),
    .Y(_01481_)
  );
  NOR2X1 _07507_ (
    .A(_01479_),
    .B(_01481_),
    .Y(_01482_)
  );
  INVX1 _07508_ (
    .A(_01482_),
    .Y(_01483_)
  );
  NAND2X1 _07509_ (
    .A(_01239_),
    .B(_01482_),
    .Y(_01484_)
  );
  AOI21X1 _07510_ (
    .A( execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01478_),
    .C(_01480_),
    .Y(_01485_)
  );
  AOI21X1 _07511_ (
    .A(_01240_),
    .B(_01481_),
    .C(_01485_),
    .Y(_01486_)
  );
  AND2X1 _07512_ (
    .A(_01484_),
    .B(_01486_),
    .Y(_01487_)
  );
  NAND2X1 _07513_ (
    .A(_01476_),
    .B(_01487_),
    .Y(_01488_)
  );
  XNOR2X1 _07514_ (
    .A(_01476_),
    .B(_01487_),
    .Y(_01489_)
  );
  INVX1 _07515_ (
    .A(_01489_),
    .Y( dbg_0.UNUSED_eu_mab_8_ )
  );
  NOR2X1 _07516_ (
    .A(_01482_),
    .B(_01485_),
    .Y(_01490_)
  );
  XNOR2X1 _07517_ (
    .A(_01416_),
    .B(_01418_),
    .Y(_01491_)
  );
  XOR2X1 _07518_ (
    .A(_01416_),
    .B(_01418_),
    .Y(_01492_)
  );
  XNOR2X1 _07519_ (
    .A(_01490_),
    .B(_01491_),
    .Y(_01493_)
  );
  AND2X1 _07520_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01490_),
    .Y(_01494_)
  );
  NAND2X1 _07521_ (
    .A(_01255_),
    .B(_01480_),
    .Y(_01495_)
  );
  AOI22X1 _07522_ (
    .A( execution_unit_0.alu_0.alu_swpb_8_ ),
    .B( execution_unit_0.alu_0.inst_so_1_ ),
    .C( execution_unit_0.alu_0.alu_shift_8_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01496_)
  );
  NAND3X1 _07523_ (
    .A(_01467_),
    .B(_01495_),
    .C(_01496_),
    .Y(_01497_)
  );
  AOI21X1 _07524_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01482_),
    .C(_01497_),
    .Y(_01498_)
  );
  OAI21X1 _07525_ (
    .A(_01219_),
    .B(_01485_),
    .C(_01498_),
    .Y(_01499_)
  );
  OAI21X1 _07526_ (
    .A(_01494_),
    .B(_01499_),
    .C(_01228_),
    .Y(_01500_)
  );
  AOI21X1 _07527_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01493_),
    .C(_01500_),
    .Y(_01501_)
  );
  INVX1 _07528_ (
    .A(_01501_),
    .Y(_01502_)
  );
  AOI21X1 _07529_ (
    .A(_01439_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .C( dbg_0.UNUSED_eu_mab_8_ ),
    .Y(_01503_)
  );
  OR2X1 _07530_ (
    .A(_01458_),
    .B(_01489_),
    .Y(_01504_)
  );
  OAI21X1 _07531_ (
    .A(_01458_),
    .B(_01489_),
    .C(_01229_),
    .Y(_01505_)
  );
  OAI21X1 _07532_ (
    .A(_01503_),
    .B(_01505_),
    .C(_01502_),
    .Y( execution_unit_0.alu_0.alu_out_8_ )
  );
  INVX1 _07533_ (
    .A( execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_01506_)
  );
  OAI21X1 _07534_ (
    .A(_01240_),
    .B(_01483_),
    .C(_01488_),
    .Y(_01507_)
  );
  XOR2X1 _07535_ (
    .A( execution_unit_0.alu_0.alu_shift_8_ ),
    .B(_01241_),
    .Y(_01508_)
  );
  NOR2X1 _07536_ (
    .A(_01477_),
    .B(_01508_),
    .Y(_01509_)
  );
  AND2X1 _07537_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01509_),
    .Y(_01510_)
  );
  NAND2X1 _07538_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01509_),
    .Y(_01511_)
  );
  NOR2X1 _07539_ (
    .A(_01240_),
    .B(_01511_),
    .Y(_01512_)
  );
  AOI21X1 _07540_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01478_),
    .C(_01509_),
    .Y(_01513_)
  );
  AOI22X1 _07541_ (
    .A( execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01478_),
    .C(_01509_),
    .D(_01239_),
    .Y(_01514_)
  );
  NOR2X1 _07542_ (
    .A(_01512_),
    .B(_01514_),
    .Y(_01515_)
  );
  XNOR2X1 _07543_ (
    .A(_01507_),
    .B(_01515_),
    .Y(_01516_)
  );
  INVX1 _07544_ (
    .A(_01516_),
    .Y( dbg_0.UNUSED_eu_mab_9_ )
  );
  AND2X1 _07545_ (
    .A(_01504_),
    .B(_01516_),
    .Y(_01517_)
  );
  OR2X1 _07546_ (
    .A(_01504_),
    .B(_01516_),
    .Y(_01518_)
  );
  OAI21X1 _07547_ (
    .A(_01504_),
    .B(_01516_),
    .C(_01229_),
    .Y(_01519_)
  );
  NOR2X1 _07548_ (
    .A(_01510_),
    .B(_01513_),
    .Y(_01520_)
  );
  AOI21X1 _07549_ (
    .A(_01490_),
    .B(_01491_),
    .C(_01482_),
    .Y(_01521_)
  );
  OAI21X1 _07550_ (
    .A(_01485_),
    .B(_01492_),
    .C(_01483_),
    .Y(_01522_)
  );
  XNOR2X1 _07551_ (
    .A(_01520_),
    .B(_01521_),
    .Y(_01523_)
  );
  XOR2X1 _07552_ (
    .A( execution_unit_0.alu_0.alu_shift_10_ ),
    .B(_01241_),
    .Y(_01524_)
  );
  NOR2X1 _07553_ (
    .A(_01477_),
    .B(_01524_),
    .Y(_01525_)
  );
  OAI21X1 _07554_ (
    .A(_01754_),
    .B(_01226_),
    .C( execution_unit_0.alu_0.op_dst_11_ ),
    .Y(_01526_)
  );
  NOR2X1 _07555_ (
    .A(_01524_),
    .B(_01526_),
    .Y(_01527_)
  );
  NAND2X1 _07556_ (
    .A( execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01525_),
    .Y(_01528_)
  );
  AOI21X1 _07557_ (
    .A( execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01478_),
    .C(_01525_),
    .Y(_01529_)
  );
  NOR2X1 _07558_ (
    .A(_01527_),
    .B(_01529_),
    .Y(_01530_)
  );
  XOR2X1 _07559_ (
    .A( execution_unit_0.alu_0.alu_shift_9_ ),
    .B(_01241_),
    .Y(_01531_)
  );
  NOR2X1 _07560_ (
    .A(_01477_),
    .B(_01531_),
    .Y(_01532_)
  );
  AND2X1 _07561_ (
    .A( execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01532_),
    .Y(_01533_)
  );
  INVX1 _07562_ (
    .A(_01533_),
    .Y(_01534_)
  );
  AOI21X1 _07563_ (
    .A( execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01478_),
    .C(_01532_),
    .Y(_01535_)
  );
  NOR2X1 _07564_ (
    .A(_01533_),
    .B(_01535_),
    .Y(_01536_)
  );
  AOI21X1 _07565_ (
    .A(_01520_),
    .B(_01522_),
    .C(_01510_),
    .Y(_01537_)
  );
  OAI21X1 _07566_ (
    .A(_01513_),
    .B(_01521_),
    .C(_01511_),
    .Y(_01538_)
  );
  AOI21X1 _07567_ (
    .A(_01536_),
    .B(_01538_),
    .C(_01533_),
    .Y(_01539_)
  );
  OAI21X1 _07568_ (
    .A(_01535_),
    .B(_01537_),
    .C(_01534_),
    .Y(_01540_)
  );
  AOI21X1 _07569_ (
    .A(_01530_),
    .B(_01540_),
    .C(_01527_),
    .Y(_01541_)
  );
  OAI21X1 _07570_ (
    .A(_01529_),
    .B(_01539_),
    .C(_01528_),
    .Y(_01542_)
  );
  XNOR2X1 _07571_ (
    .A(_01530_),
    .B(_01539_),
    .Y(_01543_)
  );
  XNOR2X1 _07572_ (
    .A(_01530_),
    .B(_01540_),
    .Y(_01544_)
  );
  XNOR2X1 _07573_ (
    .A(_01536_),
    .B(_01537_),
    .Y(_01545_)
  );
  NOR2X1 _07574_ (
    .A(_01523_),
    .B(_01545_),
    .Y(_01546_)
  );
  OR2X1 _07575_ (
    .A(_01523_),
    .B(_01545_),
    .Y(_01547_)
  );
  AOI21X1 _07576_ (
    .A(_01543_),
    .B(_01547_),
    .C(_01542_),
    .Y(_01548_)
  );
  OAI21X1 _07577_ (
    .A(_01544_),
    .B(_01546_),
    .C(_01541_),
    .Y(_01549_)
  );
  XNOR2X1 _07578_ (
    .A(_01523_),
    .B(_01548_),
    .Y(_01550_)
  );
  NAND2X1 _07579_ (
    .A(_01255_),
    .B(_01509_),
    .Y(_01551_)
  );
  AOI22X1 _07580_ (
    .A( execution_unit_0.alu_0.alu_shift_0_ ),
    .B( execution_unit_0.alu_0.inst_so_1_ ),
    .C( execution_unit_0.alu_0.alu_shift_9_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01552_)
  );
  NAND3X1 _07581_ (
    .A(_01467_),
    .B(_01551_),
    .C(_01552_),
    .Y(_01553_)
  );
  AOI21X1 _07582_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01510_),
    .C(_01553_),
    .Y(_01554_)
  );
  OAI21X1 _07583_ (
    .A(_01219_),
    .B(_01513_),
    .C(_01554_),
    .Y(_01555_)
  );
  AOI21X1 _07584_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01520_),
    .C(_01555_),
    .Y(_01556_)
  );
  NOR2X1 _07585_ (
    .A(_01229_),
    .B(_01556_),
    .Y(_01557_)
  );
  OAI21X1 _07586_ (
    .A(_01223_),
    .B(_01550_),
    .C(_01557_),
    .Y(_01558_)
  );
  OAI21X1 _07587_ (
    .A(_01517_),
    .B(_01519_),
    .C(_01558_),
    .Y( execution_unit_0.alu_0.alu_out_9_ )
  );
  INVX1 _07588_ (
    .A( execution_unit_0.alu_0.alu_out_9_ ),
    .Y(_01559_)
  );
  NOR2X1 _07589_ (
    .A(_01484_),
    .B(_01513_),
    .Y(_01560_)
  );
  NOR2X1 _07590_ (
    .A(_01512_),
    .B(_01560_),
    .Y(_01561_)
  );
  OAI21X1 _07591_ (
    .A(_01488_),
    .B(_01514_),
    .C(_01561_),
    .Y(_01562_)
  );
  AOI22X1 _07592_ (
    .A( execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01478_),
    .C(_01532_),
    .D(_01239_),
    .Y(_01563_)
  );
  AOI21X1 _07593_ (
    .A(_01239_),
    .B(_01533_),
    .C(_01563_),
    .Y(_01564_)
  );
  NAND2X1 _07594_ (
    .A(_01562_),
    .B(_01564_),
    .Y(_01565_)
  );
  XNOR2X1 _07595_ (
    .A(_01562_),
    .B(_01564_),
    .Y(_01566_)
  );
  INVX1 _07596_ (
    .A(_01566_),
    .Y( dbg_0.UNUSED_eu_mab_10_ )
  );
  NOR2X1 _07597_ (
    .A(_01518_),
    .B(_01566_),
    .Y(_01567_)
  );
  OAI21X1 _07598_ (
    .A(_01504_),
    .B(_01516_),
    .C(_01566_),
    .Y(_01568_)
  );
  OAI21X1 _07599_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01227_),
    .C(_01568_),
    .Y(_01569_)
  );
  OAI21X1 _07600_ (
    .A(_01523_),
    .B(_01548_),
    .C(_01545_),
    .Y(_01570_)
  );
  AOI21X1 _07601_ (
    .A(_01542_),
    .B(_01546_),
    .C(_01223_),
    .Y(_01571_)
  );
  NAND2X1 _07602_ (
    .A(_01570_),
    .B(_01571_),
    .Y(_01572_)
  );
  NAND2X1 _07603_ (
    .A(_01255_),
    .B(_01532_),
    .Y(_01573_)
  );
  AOI22X1 _07604_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_1_ ),
    .C( execution_unit_0.alu_0.alu_shift_10_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01574_)
  );
  NAND3X1 _07605_ (
    .A(_01467_),
    .B(_01573_),
    .C(_01574_),
    .Y(_01575_)
  );
  AOI21X1 _07606_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01533_),
    .C(_01575_),
    .Y(_01576_)
  );
  OAI21X1 _07607_ (
    .A(_01219_),
    .B(_01535_),
    .C(_01576_),
    .Y(_01577_)
  );
  AOI21X1 _07608_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01536_),
    .C(_01577_),
    .Y(_01578_)
  );
  NOR2X1 _07609_ (
    .A(_01229_),
    .B(_01578_),
    .Y(_01579_)
  );
  NAND2X1 _07610_ (
    .A(_01572_),
    .B(_01579_),
    .Y(_01580_)
  );
  OAI21X1 _07611_ (
    .A(_01567_),
    .B(_01569_),
    .C(_01580_),
    .Y( execution_unit_0.alu_0.alu_out_10_ )
  );
  NAND2X1 _07612_ (
    .A(_01239_),
    .B(_01525_),
    .Y(_01581_)
  );
  AOI22X1 _07613_ (
    .A(_01239_),
    .B(_01527_),
    .C(_01581_),
    .D(_01526_),
    .Y(_01582_)
  );
  OAI21X1 _07614_ (
    .A(_01240_),
    .B(_01534_),
    .C(_01565_),
    .Y(_01583_)
  );
  NAND2X1 _07615_ (
    .A(_01582_),
    .B(_01583_),
    .Y(_01584_)
  );
  XOR2X1 _07616_ (
    .A(_01582_),
    .B(_01583_),
    .Y( dbg_0.UNUSED_eu_mab_11_ )
  );
  NAND2X1 _07617_ (
    .A(_01567_),
    .B( dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_01585_)
  );
  XOR2X1 _07618_ (
    .A(_01567_),
    .B( dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_01586_)
  );
  AOI22X1 _07619_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.alu_shift_11_ ),
    .C( execution_unit_0.alu_0.alu_shift_6_ ),
    .D( execution_unit_0.alu_0.inst_so_3_ ),
    .Y(_01587_)
  );
  AOI22X1 _07620_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_2_ ),
    .C(_01255_),
    .D(_01525_),
    .Y(_01588_)
  );
  OAI21X1 _07621_ (
    .A(_01218_),
    .B(_01528_),
    .C(_01588_),
    .Y(_01589_)
  );
  OAI21X1 _07622_ (
    .A(_01219_),
    .B(_01529_),
    .C(_01587_),
    .Y(_01590_)
  );
  NOR2X1 _07623_ (
    .A(_01589_),
    .B(_01590_),
    .Y(_01591_)
  );
  AOI21X1 _07624_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01530_),
    .C(_01229_),
    .Y(_01592_)
  );
  AOI22X1 _07625_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01228_),
    .C(_01591_),
    .D(_01592_),
    .Y(_01593_)
  );
  AOI21X1 _07626_ (
    .A(_01542_),
    .B(_01547_),
    .C(_01543_),
    .Y(_01594_)
  );
  OAI21X1 _07627_ (
    .A(_01544_),
    .B(_01546_),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01595_)
  );
  NOR2X1 _07628_ (
    .A(_01594_),
    .B(_01595_),
    .Y(_01596_)
  );
  OAI22X1 _07629_ (
    .A(_01228_),
    .B(_01586_),
    .C(_01593_),
    .D(_01596_),
    .Y(_01597_)
  );
  INVX1 _07630_ (
    .A(_01597_),
    .Y( execution_unit_0.alu_0.alu_out_11_ )
  );
  OAI21X1 _07631_ (
    .A(_01240_),
    .B(_01528_),
    .C(_01584_),
    .Y(_01598_)
  );
  XOR2X1 _07632_ (
    .A( execution_unit_0.alu_0.alu_shift_11_ ),
    .B(_01241_),
    .Y(_01599_)
  );
  NOR2X1 _07633_ (
    .A(_01477_),
    .B(_01599_),
    .Y(_01600_)
  );
  AND2X1 _07634_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01600_),
    .Y(_01601_)
  );
  NAND2X1 _07635_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01600_),
    .Y(_01602_)
  );
  NAND2X1 _07636_ (
    .A(_01239_),
    .B(_01601_),
    .Y(_01603_)
  );
  AOI21X1 _07637_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01478_),
    .C(_01600_),
    .Y(_01604_)
  );
  AOI22X1 _07638_ (
    .A( execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01478_),
    .C(_01600_),
    .D(_01239_),
    .Y(_01605_)
  );
  AOI21X1 _07639_ (
    .A(_01239_),
    .B(_01601_),
    .C(_01605_),
    .Y(_01606_)
  );
  NAND2X1 _07640_ (
    .A(_01598_),
    .B(_01606_),
    .Y(_01607_)
  );
  XNOR2X1 _07641_ (
    .A(_01598_),
    .B(_01606_),
    .Y(_01608_)
  );
  INVX1 _07642_ (
    .A(_01608_),
    .Y( dbg_0.UNUSED_eu_mab_12_ )
  );
  NOR2X1 _07643_ (
    .A(_01585_),
    .B(_01608_),
    .Y(_01609_)
  );
  NAND2X1 _07644_ (
    .A(_01585_),
    .B(_01608_),
    .Y(_01610_)
  );
  OAI21X1 _07645_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01227_),
    .C(_01610_),
    .Y(_01611_)
  );
  NOR2X1 _07646_ (
    .A(_01601_),
    .B(_01604_),
    .Y(_01612_)
  );
  INVX1 _07647_ (
    .A(_01612_),
    .Y(_01613_)
  );
  NOR3X1 _07648_ (
    .A(_01541_),
    .B(_01544_),
    .C(_01546_),
    .Y(_01614_)
  );
  NAND3X1 _07649_ (
    .A(_01542_),
    .B(_01543_),
    .C(_01547_),
    .Y(_01615_)
  );
  OAI21X1 _07650_ (
    .A(_01548_),
    .B(_01614_),
    .C(_01613_),
    .Y(_01616_)
  );
  NOR3X1 _07651_ (
    .A(_01548_),
    .B(_01613_),
    .C(_01614_),
    .Y(_01617_)
  );
  NAND3X1 _07652_ (
    .A(_01549_),
    .B(_01612_),
    .C(_01615_),
    .Y(_01618_)
  );
  AND2X1 _07653_ (
    .A(_01616_),
    .B(_01618_),
    .Y(_01619_)
  );
  NAND2X1 _07654_ (
    .A(_01255_),
    .B(_01600_),
    .Y(_01620_)
  );
  AOI22X1 _07655_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_3_ ),
    .C( execution_unit_0.alu_0.alu_shift_12_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01621_)
  );
  NAND3X1 _07656_ (
    .A(_01467_),
    .B(_01620_),
    .C(_01621_),
    .Y(_01622_)
  );
  AOI21X1 _07657_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01601_),
    .C(_01622_),
    .Y(_01623_)
  );
  OAI21X1 _07658_ (
    .A(_01219_),
    .B(_01604_),
    .C(_01623_),
    .Y(_01624_)
  );
  AOI21X1 _07659_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01612_),
    .C(_01624_),
    .Y(_01625_)
  );
  NOR2X1 _07660_ (
    .A(_01229_),
    .B(_01625_),
    .Y(_01626_)
  );
  OAI21X1 _07661_ (
    .A(_01223_),
    .B(_01619_),
    .C(_01626_),
    .Y(_01627_)
  );
  OAI21X1 _07662_ (
    .A(_01609_),
    .B(_01611_),
    .C(_01627_),
    .Y( execution_unit_0.alu_0.alu_out_12_ )
  );
  OAI21X1 _07663_ (
    .A(_01240_),
    .B(_01602_),
    .C(_01607_),
    .Y(_01628_)
  );
  XOR2X1 _07664_ (
    .A( execution_unit_0.alu_0.alu_shift_12_ ),
    .B(_01241_),
    .Y(_01629_)
  );
  NOR2X1 _07665_ (
    .A(_01477_),
    .B(_01629_),
    .Y(_01630_)
  );
  AND2X1 _07666_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01630_),
    .Y(_01631_)
  );
  NAND2X1 _07667_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01630_),
    .Y(_01632_)
  );
  AOI21X1 _07668_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01478_),
    .C(_01630_),
    .Y(_01633_)
  );
  AOI22X1 _07669_ (
    .A( execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01478_),
    .C(_01630_),
    .D(_01239_),
    .Y(_01634_)
  );
  AOI21X1 _07670_ (
    .A(_01239_),
    .B(_01631_),
    .C(_01634_),
    .Y(_01635_)
  );
  XOR2X1 _07671_ (
    .A(_01628_),
    .B(_01635_),
    .Y( dbg_0.UNUSED_eu_mab_13_ )
  );
  AND2X1 _07672_ (
    .A(_01609_),
    .B( dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01636_)
  );
  XNOR2X1 _07673_ (
    .A(_01609_),
    .B( dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01637_)
  );
  NOR2X1 _07674_ (
    .A(_01631_),
    .B(_01633_),
    .Y(_01638_)
  );
  INVX1 _07675_ (
    .A(_01638_),
    .Y(_01639_)
  );
  NAND2X1 _07676_ (
    .A(_01602_),
    .B(_01618_),
    .Y(_01640_)
  );
  AOI21X1 _07677_ (
    .A(_01602_),
    .B(_01618_),
    .C(_01639_),
    .Y(_01641_)
  );
  OAI21X1 _07678_ (
    .A(_01601_),
    .B(_01617_),
    .C(_01638_),
    .Y(_01642_)
  );
  XNOR2X1 _07679_ (
    .A(_01639_),
    .B(_01640_),
    .Y(_01643_)
  );
  XNOR2X1 _07680_ (
    .A(_01638_),
    .B(_01640_),
    .Y(_01644_)
  );
  XOR2X1 _07681_ (
    .A( execution_unit_0.alu_0.alu_shift_14_ ),
    .B(_01241_),
    .Y(_01645_)
  );
  NOR2X1 _07682_ (
    .A(_01477_),
    .B(_01645_),
    .Y(_01646_)
  );
  OAI21X1 _07683_ (
    .A(_01754_),
    .B(_01226_),
    .C( execution_unit_0.alu_0.op_dst_15_ ),
    .Y(_01647_)
  );
  NOR2X1 _07684_ (
    .A(_01645_),
    .B(_01647_),
    .Y(_01648_)
  );
  NAND2X1 _07685_ (
    .A( execution_unit_0.alu_0.op_dst_15_ ),
    .B(_01646_),
    .Y(_01649_)
  );
  OAI21X1 _07686_ (
    .A(_01477_),
    .B(_01645_),
    .C(_01647_),
    .Y(_01650_)
  );
  XOR2X1 _07687_ (
    .A( execution_unit_0.alu_0.alu_shift_13_ ),
    .B(_01241_),
    .Y(_01651_)
  );
  NOR2X1 _07688_ (
    .A(_01477_),
    .B(_01651_),
    .Y(_01652_)
  );
  AND2X1 _07689_ (
    .A( execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01478_),
    .Y(_01653_)
  );
  AND2X1 _07690_ (
    .A( execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01652_),
    .Y(_01654_)
  );
  NAND2X1 _07691_ (
    .A( execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01652_),
    .Y(_01655_)
  );
  NOR2X1 _07692_ (
    .A(_01652_),
    .B(_01653_),
    .Y(_01656_)
  );
  NOR2X1 _07693_ (
    .A(_01654_),
    .B(_01656_),
    .Y(_01657_)
  );
  OAI21X1 _07694_ (
    .A(_01652_),
    .B(_01653_),
    .C(_01655_),
    .Y(_01658_)
  );
  AOI21X1 _07695_ (
    .A(_01632_),
    .B(_01642_),
    .C(_01658_),
    .Y(_01659_)
  );
  OAI21X1 _07696_ (
    .A(_01631_),
    .B(_01641_),
    .C(_01657_),
    .Y(_01660_)
  );
  OAI21X1 _07697_ (
    .A(_01654_),
    .B(_01659_),
    .C(_01650_),
    .Y(_01661_)
  );
  AND2X1 _07698_ (
    .A(_01649_),
    .B(_01661_),
    .Y(_01662_)
  );
  OAI21X1 _07699_ (
    .A(_01645_),
    .B(_01647_),
    .C(_01661_),
    .Y(_01663_)
  );
  NOR3X1 _07700_ (
    .A(_01631_),
    .B(_01641_),
    .C(_01657_),
    .Y(_01664_)
  );
  NAND3X1 _07701_ (
    .A(_01632_),
    .B(_01642_),
    .C(_01658_),
    .Y(_01665_)
  );
  NOR2X1 _07702_ (
    .A(_01659_),
    .B(_01664_),
    .Y(_01666_)
  );
  AOI21X1 _07703_ (
    .A(_01660_),
    .B(_01665_),
    .C(_01643_),
    .Y(_01667_)
  );
  OAI21X1 _07704_ (
    .A(_01659_),
    .B(_01664_),
    .C(_01644_),
    .Y(_01668_)
  );
  AND2X1 _07705_ (
    .A(_01649_),
    .B(_01650_),
    .Y(_01669_)
  );
  OAI21X1 _07706_ (
    .A(_01645_),
    .B(_01647_),
    .C(_01650_),
    .Y(_01670_)
  );
  NOR3X1 _07707_ (
    .A(_01654_),
    .B(_01659_),
    .C(_01669_),
    .Y(_01671_)
  );
  NAND3X1 _07708_ (
    .A(_01655_),
    .B(_01660_),
    .C(_01670_),
    .Y(_01672_)
  );
  AOI21X1 _07709_ (
    .A(_01655_),
    .B(_01660_),
    .C(_01670_),
    .Y(_01673_)
  );
  OAI21X1 _07710_ (
    .A(_01654_),
    .B(_01659_),
    .C(_01669_),
    .Y(_01674_)
  );
  NOR3X1 _07711_ (
    .A(_01667_),
    .B(_01671_),
    .C(_01673_),
    .Y(_01675_)
  );
  NAND3X1 _07712_ (
    .A(_01668_),
    .B(_01672_),
    .C(_01674_),
    .Y(_01676_)
  );
  AOI21X1 _07713_ (
    .A(_01662_),
    .B(_01676_),
    .C(_01643_),
    .Y(_01677_)
  );
  OAI21X1 _07714_ (
    .A(_01663_),
    .B(_01675_),
    .C(_01644_),
    .Y(_01678_)
  );
  NOR3X1 _07715_ (
    .A(_01644_),
    .B(_01663_),
    .C(_01675_),
    .Y(_01679_)
  );
  NOR3X1 _07716_ (
    .A(_01223_),
    .B(_01677_),
    .C(_01679_),
    .Y(_01680_)
  );
  NOR2X1 _07717_ (
    .A(_01220_),
    .B(_01639_),
    .Y(_01681_)
  );
  NAND2X1 _07718_ (
    .A(_01255_),
    .B(_01630_),
    .Y(_01682_)
  );
  AOI22X1 _07719_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_4_ ),
    .C( execution_unit_0.alu_0.alu_shift_13_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01683_)
  );
  NAND3X1 _07720_ (
    .A(_01467_),
    .B(_01682_),
    .C(_01683_),
    .Y(_01684_)
  );
  AOI21X1 _07721_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01631_),
    .C(_01684_),
    .Y(_01685_)
  );
  OAI21X1 _07722_ (
    .A(_01219_),
    .B(_01633_),
    .C(_01685_),
    .Y(_01686_)
  );
  OAI21X1 _07723_ (
    .A(_01681_),
    .B(_01686_),
    .C(_01228_),
    .Y(_01687_)
  );
  OAI22X1 _07724_ (
    .A(_01228_),
    .B(_01637_),
    .C(_01680_),
    .D(_01687_),
    .Y( execution_unit_0.alu_0.alu_out_13_ )
  );
  OAI22X1 _07725_ (
    .A(_01240_),
    .B(_01632_),
    .C(_01633_),
    .D(_01603_),
    .Y(_01688_)
  );
  INVX1 _07726_ (
    .A(_01688_),
    .Y(_01689_)
  );
  OAI21X1 _07727_ (
    .A(_01607_),
    .B(_01634_),
    .C(_01689_),
    .Y(_01690_)
  );
  AOI21X1 _07728_ (
    .A(_01239_),
    .B(_01652_),
    .C(_01653_),
    .Y(_01691_)
  );
  AOI21X1 _07729_ (
    .A(_01239_),
    .B(_01654_),
    .C(_01691_),
    .Y(_01692_)
  );
  NAND2X1 _07730_ (
    .A(_01690_),
    .B(_01692_),
    .Y(_01693_)
  );
  XOR2X1 _07731_ (
    .A(_01690_),
    .B(_01692_),
    .Y( dbg_0.UNUSED_eu_mab_14_ )
  );
  OAI21X1 _07732_ (
    .A(_01662_),
    .B(_01668_),
    .C( execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01694_)
  );
  AOI21X1 _07733_ (
    .A(_01666_),
    .B(_01678_),
    .C(_01694_),
    .Y(_01695_)
  );
  OAI21X1 _07734_ (
    .A(_01652_),
    .B(_01653_),
    .C( execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01696_)
  );
  AOI22X1 _07735_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B( execution_unit_0.alu_0.alu_shift_6_ ),
    .C( execution_unit_0.alu_0.alu_shift_14_ ),
    .D( execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01697_)
  );
  AOI22X1 _07736_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.alu_shift_5_ ),
    .C(_01255_),
    .D(_01652_),
    .Y(_01698_)
  );
  OAI21X1 _07737_ (
    .A(_01218_),
    .B(_01655_),
    .C(_01698_),
    .Y(_01699_)
  );
  AOI21X1 _07738_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01657_),
    .C(_01699_),
    .Y(_01700_)
  );
  NAND3X1 _07739_ (
    .A(_01696_),
    .B(_01697_),
    .C(_01700_),
    .Y(_01701_)
  );
  OAI21X1 _07740_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01701_),
    .C(_01228_),
    .Y(_01702_)
  );
  AND2X1 _07741_ (
    .A(_01636_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .Y(_01703_)
  );
  NAND2X1 _07742_ (
    .A(_01636_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .Y(_01704_)
  );
  OAI21X1 _07743_ (
    .A(_01636_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .C(_01229_),
    .Y(_01705_)
  );
  OAI22X1 _07744_ (
    .A(_01695_),
    .B(_01702_),
    .C(_01703_),
    .D(_01705_),
    .Y( execution_unit_0.alu_0.alu_out_14_ )
  );
  NAND2X1 _07745_ (
    .A(_01239_),
    .B(_01646_),
    .Y(_01706_)
  );
  AOI22X1 _07746_ (
    .A(_01239_),
    .B(_01648_),
    .C(_01706_),
    .D(_01647_),
    .Y(_01707_)
  );
  OAI21X1 _07747_ (
    .A(_01240_),
    .B(_01655_),
    .C(_01693_),
    .Y(_01708_)
  );
  XOR2X1 _07748_ (
    .A(_01707_),
    .B(_01708_),
    .Y( dbg_0.UNUSED_eu_mab_15_ )
  );
  INVX1 _07749_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_01709_)
  );
  XNOR2X1 _07750_ (
    .A(_01704_),
    .B( dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_01710_)
  );
  NOR2X1 _07751_ (
    .A(_01228_),
    .B(_01710_),
    .Y(_01711_)
  );
  AND2X1 _07752_ (
    .A(_01255_),
    .B(_01646_),
    .Y(_01712_)
  );
  OAI21X1 _07753_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B( execution_unit_0.alu_0.inst_so_3_ ),
    .C( execution_unit_0.alu_0.alu_shift_6_ ),
    .Y(_01713_)
  );
  OAI21X1 _07754_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01712_),
    .C(_01650_),
    .Y(_01714_)
  );
  OAI22X1 _07755_ (
    .A(_01221_),
    .B(_01464_),
    .C(_01649_),
    .D(_01218_),
    .Y(_01715_)
  );
  AOI21X1 _07756_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01669_),
    .C(_01715_),
    .Y(_01716_)
  );
  NAND3X1 _07757_ (
    .A(_01713_),
    .B(_01714_),
    .C(_01716_),
    .Y(_01717_)
  );
  INVX1 _07758_ (
    .A(_01717_),
    .Y(_01718_)
  );
  OAI21X1 _07759_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01718_),
    .C(_01228_),
    .Y(_01719_)
  );
  OAI22X1 _07760_ (
    .A(_01662_),
    .B(_01667_),
    .C(_01671_),
    .D(_01673_),
    .Y(_01720_)
  );
  NOR2X1 _07761_ (
    .A(_01223_),
    .B(_01675_),
    .Y(_01721_)
  );
  AOI21X1 _07762_ (
    .A(_01720_),
    .B(_01721_),
    .C(_01719_),
    .Y(_01722_)
  );
  NOR2X1 _07763_ (
    .A(_01711_),
    .B(_01722_),
    .Y( execution_unit_0.alu_0.alu_out_15_ )
  );
  NAND2X1 _07764_ (
    .A(_01226_),
    .B( execution_unit_0.alu_0.alu_out_15_ ),
    .Y(_01723_)
  );
  OAI21X1 _07765_ (
    .A(_01226_),
    .B(_01474_),
    .C(_01723_),
    .Y( execution_unit_0.alu_0.N )
  );
  NAND3X1 _07766_ (
    .A(_01506_),
    .B(_01559_),
    .C(_01597_),
    .Y(_01724_)
  );
  OR2X1 _07767_ (
    .A( execution_unit_0.alu_0.alu_out_10_ ),
    .B(_01724_),
    .Y(_01725_)
  );
  NOR2X1 _07768_ (
    .A( execution_unit_0.alu_0.alu_out_12_ ),
    .B(_01725_),
    .Y(_01726_)
  );
  OAI21X1 _07769_ (
    .A(_01711_),
    .B(_01722_),
    .C(_01726_),
    .Y(_01727_)
  );
  NOR3X1 _07770_ (
    .A( execution_unit_0.alu_0.alu_out_13_ ),
    .B( execution_unit_0.alu_0.alu_out_14_ ),
    .C(_01727_),
    .Y(_01728_)
  );
  OR2X1 _07771_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_01729_)
  );
  NOR2X1 _07772_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_01729_),
    .Y(_01730_)
  );
  NOR2X1 _07773_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_01731_)
  );
  NAND3X1 _07774_ (
    .A(_01474_),
    .B(_01730_),
    .C(_01731_),
    .Y(_01732_)
  );
  NOR3X1 _07775_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B( execution_unit_0.alu_0.alu_out_6_ ),
    .C(_01732_),
    .Y(_01733_)
  );
  OAI21X1 _07776_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_01728_),
    .C(_01733_),
    .Y(_01734_)
  );
  INVX1 _07777_ (
    .A(_01734_),
    .Y( execution_unit_0.alu_0.Z )
  );
  NAND2X1 _07778_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_01242_),
    .Y(_01735_)
  );
  NOR2X1 _07779_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B( execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01736_)
  );
  NOR2X1 _07780_ (
    .A(_01734_),
    .B(_01736_),
    .Y(_01737_)
  );
  AOI22X1 _07781_ (
    .A(_01239_),
    .B(_01648_),
    .C(_01707_),
    .D(_01708_),
    .Y(_01738_)
  );
  OAI21X1 _07782_ (
    .A(_01704_),
    .B(_01709_),
    .C(_01738_),
    .Y(_01739_)
  );
  OAI21X1 _07783_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01227_),
    .C(_01739_),
    .Y(_01740_)
  );
  AOI21X1 _07784_ (
    .A(_01662_),
    .B(_01676_),
    .C(_01324_),
    .Y(_01741_)
  );
  OAI21X1 _07785_ (
    .A(_01662_),
    .B(_01676_),
    .C(_01741_),
    .Y(_01742_)
  );
  AOI21X1 _07786_ (
    .A(_01740_),
    .B(_01742_),
    .C( execution_unit_0.alu_0.inst_bw ),
    .Y(_01743_)
  );
  OAI21X1 _07787_ (
    .A(_01226_),
    .B(_01506_),
    .C(_01736_),
    .Y(_01744_)
  );
  OAI21X1 _07788_ (
    .A(_01743_),
    .B(_01744_),
    .C(_01221_),
    .Y(_01745_)
  );
  OAI21X1 _07789_ (
    .A(_01737_),
    .B(_01745_),
    .C(_01735_),
    .Y( execution_unit_0.alu_0.alu_stat_0_ )
  );
  NOR2X1 _07790_ (
    .A(_01409_),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01746_)
  );
  OAI21X1 _07791_ (
    .A(_01410_),
    .B(_01474_),
    .C( execution_unit_0.alu_0.inst_bw ),
    .Y(_01747_)
  );
  MUX2X1 _07792_ (
    .A(_01650_),
    .B(_01649_),
    .S( execution_unit_0.alu_0.alu_out_15_ ),
    .Y(_01748_)
  );
  OAI22X1 _07793_ (
    .A(_01746_),
    .B(_01747_),
    .C(_01748_),
    .D( execution_unit_0.alu_0.inst_bw ),
    .Y(_01749_)
  );
  NOR2X1 _07794_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_01649_),
    .Y(_01750_)
  );
  OAI21X1 _07795_ (
    .A(_01226_),
    .B(_01409_),
    .C( execution_unit_0.alu_0.inst_alu_6_ ),
    .Y(_01751_)
  );
  NOR2X1 _07796_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B( execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01752_)
  );
  OAI21X1 _07797_ (
    .A(_01750_),
    .B(_01751_),
    .C(_01752_),
    .Y(_01753_)
  );
  AOI21X1 _07798_ (
    .A(_01220_),
    .B(_01749_),
    .C(_01753_),
    .Y( execution_unit_0.alu_0.alu_stat_3_ )
  );
  AND2X1 _07799_ (
    .A( execution_unit_0.alu_0.exec_cycle ),
    .B( execution_unit_0.alu_0.inst_alu_9_ ),
    .Y( execution_unit_0.alu_0.alu_stat_wr_0_ )
  );
  INVX1 _07800_ (
    .A( execution_unit_0.reg_sp_wr ),
    .Y(_02539_)
  );
  INVX1 _07801_ (
    .A( execution_unit_0.reg_sr_clr ),
    .Y(_02540_)
  );
  INVX1 _07802_ (
    .A( execution_unit_0.inst_src_1_ ),
    .Y(_02541_)
  );
  INVX1 _07803_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_02542_)
  );
  INVX1 _07804_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_02543_)
  );
  INVX1 _07805_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .Y(_02544_)
  );
  INVX1 _07806_ (
    .A( execution_unit_0.register_file_0.r5_0_ ),
    .Y(_02545_)
  );
  INVX1 _07807_ (
    .A( execution_unit_0.register_file_0.r6_0_ ),
    .Y(_02546_)
  );
  INVX1 _07808_ (
    .A( execution_unit_0.register_file_0.r7_0_ ),
    .Y(_02547_)
  );
  INVX1 _07809_ (
    .A( execution_unit_0.register_file_0.r8_0_ ),
    .Y(_02548_)
  );
  INVX1 _07810_ (
    .A( execution_unit_0.register_file_0.r10_0_ ),
    .Y(_02549_)
  );
  INVX1 _07811_ (
    .A( execution_unit_0.register_file_0.r11_0_ ),
    .Y(_02550_)
  );
  INVX1 _07812_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_02551_)
  );
  INVX1 _07813_ (
    .A( execution_unit_0.register_file_0.r6_1_ ),
    .Y(_02552_)
  );
  INVX1 _07814_ (
    .A( execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02553_)
  );
  INVX1 _07815_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_02554_)
  );
  INVX1 _07816_ (
    .A( execution_unit_0.register_file_0.r10_2_ ),
    .Y(_02555_)
  );
  INVX1 _07817_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_02556_)
  );
  INVX1 _07818_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_02557_)
  );
  INVX1 _07819_ (
    .A( execution_unit_0.register_file_0.r2_4_ ),
    .Y(_02558_)
  );
  INVX1 _07820_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_02559_)
  );
  INVX1 _07821_ (
    .A( execution_unit_0.register_file_0.r11_5_ ),
    .Y(_02560_)
  );
  INVX1 _07822_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_02561_)
  );
  INVX1 _07823_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .Y(_02562_)
  );
  INVX1 _07824_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_02563_)
  );
  INVX1 _07825_ (
    .A( execution_unit_0.register_file_0.r6_15_ ),
    .Y(_02564_)
  );
  INVX1 _07826_ (
    .A(_05695_),
    .Y(_01756_)
  );
  OR2X1 _07827_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .Y(_02565_)
  );
  NOR2X1 _07828_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B(_02541_),
    .Y(_02566_)
  );
  AOI22X1 _07829_ (
    .A( execution_unit_0.gie ),
    .B(_02565_),
    .C(_02566_),
    .D( execution_unit_0.register_file_0.r1_3_ ),
    .Y(_02567_)
  );
  AND2X1 _07830_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_13_ ),
    .Y(_02568_)
  );
  AND2X1 _07831_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_15_ ),
    .Y(_02569_)
  );
  AOI22X1 _07832_ (
    .A( execution_unit_0.register_file_0.r13_3_ ),
    .B(_02568_),
    .C(_02569_),
    .D( execution_unit_0.register_file_0.r15_3_ ),
    .Y(_02570_)
  );
  AND2X1 _07833_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_4_ ),
    .Y(_02571_)
  );
  AND2X1 _07834_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_0_ ),
    .Y(_02572_)
  );
  AOI22X1 _07835_ (
    .A( execution_unit_0.register_file_0.r4_3_ ),
    .B(_02571_),
    .C(_02572_),
    .D( dbg_0.UNUSED_pc_3_ ),
    .Y(_02573_)
  );
  AND2X1 _07836_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_3_ ),
    .Y(_02574_)
  );
  AND2X1 _07837_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_6_ ),
    .Y(_02575_)
  );
  NAND2X1 _07838_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_6_ ),
    .Y(_02576_)
  );
  AOI22X1 _07839_ (
    .A( execution_unit_0.register_file_0.r3_3_ ),
    .B(_02574_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_3_ ),
    .Y(_02577_)
  );
  AND2X1 _07840_ (
    .A(_02573_),
    .B(_02577_),
    .Y(_02578_)
  );
  NAND3X1 _07841_ (
    .A(_02567_),
    .B(_02570_),
    .C(_02578_),
    .Y(_02579_)
  );
  AND2X1 _07842_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_14_ ),
    .Y(_02580_)
  );
  AND2X1 _07843_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_8_ ),
    .Y(_02581_)
  );
  AOI22X1 _07844_ (
    .A( execution_unit_0.register_file_0.r14_3_ ),
    .B(_02580_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_3_ ),
    .Y(_02582_)
  );
  AND2X1 _07845_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_10_ ),
    .Y(_02583_)
  );
  NAND2X1 _07846_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_10_ ),
    .Y(_02584_)
  );
  AND2X1 _07847_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_7_ ),
    .Y(_02585_)
  );
  NAND2X1 _07848_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_7_ ),
    .Y(_02586_)
  );
  AOI22X1 _07849_ (
    .A( execution_unit_0.register_file_0.r10_3_ ),
    .B(_02583_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02587_)
  );
  AND2X1 _07850_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_9_ ),
    .Y(_02588_)
  );
  AND2X1 _07851_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_5_ ),
    .Y(_02589_)
  );
  AOI22X1 _07852_ (
    .A( execution_unit_0.register_file_0.r9_3_ ),
    .B(_02588_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_3_ ),
    .Y(_02590_)
  );
  AND2X1 _07853_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_11_ ),
    .Y(_02591_)
  );
  NAND2X1 _07854_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_11_ ),
    .Y(_02592_)
  );
  AND2X1 _07855_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_12_ ),
    .Y(_02593_)
  );
  AOI22X1 _07856_ (
    .A( execution_unit_0.register_file_0.r11_3_ ),
    .B(_02591_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_3_ ),
    .Y(_02594_)
  );
  AND2X1 _07857_ (
    .A(_02590_),
    .B(_02594_),
    .Y(_02595_)
  );
  NAND3X1 _07858_ (
    .A(_02582_),
    .B(_02587_),
    .C(_02595_),
    .Y(_02596_)
  );
  NOR2X1 _07859_ (
    .A(_02579_),
    .B(_02596_),
    .Y(_02597_)
  );
  INVX1 _07860_ (
    .A(_02597_),
    .Y( execution_unit_0.reg_src_3_ )
  );
  NAND2X1 _07861_ (
    .A( execution_unit_0.register_file_0.r5_2_ ),
    .B(_02589_),
    .Y(_02598_)
  );
  NAND2X1 _07862_ (
    .A( execution_unit_0.register_file_0.r13_2_ ),
    .B(_02568_),
    .Y(_02599_)
  );
  OAI21X1 _07863_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .C( execution_unit_0.alu_0.status_2_ ),
    .Y(_02600_)
  );
  AOI22X1 _07864_ (
    .A( execution_unit_0.register_file_0.r3_2_ ),
    .B(_02574_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_2_ ),
    .Y(_02601_)
  );
  NAND3X1 _07865_ (
    .A(_02598_),
    .B(_02600_),
    .C(_02601_),
    .Y(_02602_)
  );
  AOI22X1 _07866_ (
    .A( execution_unit_0.register_file_0.r4_2_ ),
    .B(_02571_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_2_ ),
    .Y(_02603_)
  );
  AOI22X1 _07867_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .B(_02572_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_2_ ),
    .Y(_02604_)
  );
  NAND2X1 _07868_ (
    .A(_02603_),
    .B(_02604_),
    .Y(_02605_)
  );
  NOR2X1 _07869_ (
    .A(_02602_),
    .B(_02605_),
    .Y(_02606_)
  );
  AOI22X1 _07870_ (
    .A( execution_unit_0.register_file_0.r11_2_ ),
    .B(_02591_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_2_ ),
    .Y(_02607_)
  );
  OAI21X1 _07871_ (
    .A(_02555_),
    .B(_02584_),
    .C(_02607_),
    .Y(_02608_)
  );
  AOI22X1 _07872_ (
    .A( execution_unit_0.register_file_0.r14_2_ ),
    .B(_02580_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_2_ ),
    .Y(_02609_)
  );
  AOI22X1 _07873_ (
    .A( execution_unit_0.register_file_0.r1_2_ ),
    .B(_02566_),
    .C(_02569_),
    .D( execution_unit_0.register_file_0.r15_2_ ),
    .Y(_02610_)
  );
  NAND3X1 _07874_ (
    .A(_02599_),
    .B(_02609_),
    .C(_02610_),
    .Y(_02611_)
  );
  NOR2X1 _07875_ (
    .A(_02608_),
    .B(_02611_),
    .Y(_02612_)
  );
  AND2X1 _07876_ (
    .A(_02606_),
    .B(_02612_),
    .Y(_02613_)
  );
  INVX1 _07877_ (
    .A(_02613_),
    .Y( execution_unit_0.reg_src_2_ )
  );
  OAI21X1 _07878_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .C( execution_unit_0.register_file_0.r2_4_ ),
    .Y(_02614_)
  );
  AOI22X1 _07879_ (
    .A( execution_unit_0.register_file_0.r10_4_ ),
    .B(_02583_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_4_ ),
    .Y(_02615_)
  );
  AOI22X1 _07880_ (
    .A( execution_unit_0.register_file_0.r15_4_ ),
    .B(_02569_),
    .C(_02574_),
    .D( execution_unit_0.register_file_0.r3_4_ ),
    .Y(_02616_)
  );
  AOI22X1 _07881_ (
    .A( execution_unit_0.register_file_0.r13_4_ ),
    .B(_02568_),
    .C(_02580_),
    .D( execution_unit_0.register_file_0.r14_4_ ),
    .Y(_02617_)
  );
  NAND2X1 _07882_ (
    .A(_02614_),
    .B(_02617_),
    .Y(_02618_)
  );
  AOI22X1 _07883_ (
    .A( execution_unit_0.register_file_0.r4_4_ ),
    .B(_02571_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_4_ ),
    .Y(_02619_)
  );
  AOI22X1 _07884_ (
    .A( execution_unit_0.register_file_0.r8_4_ ),
    .B(_02581_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_4_ ),
    .Y(_02620_)
  );
  NAND2X1 _07885_ (
    .A(_02619_),
    .B(_02620_),
    .Y(_02621_)
  );
  AOI22X1 _07886_ (
    .A( execution_unit_0.register_file_0.r1_4_ ),
    .B(_02566_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_4_ ),
    .Y(_02622_)
  );
  NAND2X1 _07887_ (
    .A(_02615_),
    .B(_02622_),
    .Y(_02623_)
  );
  NOR2X1 _07888_ (
    .A(_02621_),
    .B(_02623_),
    .Y(_02624_)
  );
  AOI22X1 _07889_ (
    .A( execution_unit_0.register_file_0.r9_4_ ),
    .B(_02588_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_4_ ),
    .Y(_02625_)
  );
  NAND2X1 _07890_ (
    .A(_02616_),
    .B(_02625_),
    .Y(_02626_)
  );
  AOI21X1 _07891_ (
    .A( dbg_0.UNUSED_pc_4_ ),
    .B(_02572_),
    .C(_02626_),
    .Y(_02627_)
  );
  NAND2X1 _07892_ (
    .A(_02624_),
    .B(_02627_),
    .Y(_02628_)
  );
  NOR2X1 _07893_ (
    .A(_02618_),
    .B(_02628_),
    .Y(_02629_)
  );
  INVX1 _07894_ (
    .A(_02629_),
    .Y( execution_unit_0.reg_src_4_ )
  );
  NAND2X1 _07895_ (
    .A( execution_unit_0.register_file_0.r13_5_ ),
    .B(_02568_),
    .Y(_02630_)
  );
  NAND2X1 _07896_ (
    .A( dbg_0.UNUSED_pc_5_ ),
    .B(_02572_),
    .Y(_02631_)
  );
  NAND2X1 _07897_ (
    .A( execution_unit_0.register_file_0.r12_5_ ),
    .B(_02593_),
    .Y(_02632_)
  );
  AOI22X1 _07898_ (
    .A( execution_unit_0.register_file_0.r15_5_ ),
    .B(_02569_),
    .C(_02580_),
    .D( execution_unit_0.register_file_0.r14_5_ ),
    .Y(_02633_)
  );
  AOI22X1 _07899_ (
    .A( clock_module_0.oscoff ),
    .B(_02565_),
    .C(_02571_),
    .D( execution_unit_0.register_file_0.r4_5_ ),
    .Y(_02634_)
  );
  AOI22X1 _07900_ (
    .A( execution_unit_0.register_file_0.r3_5_ ),
    .B(_02574_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_5_ ),
    .Y(_02635_)
  );
  NAND2X1 _07901_ (
    .A(_02634_),
    .B(_02635_),
    .Y(_02636_)
  );
  AOI21X1 _07902_ (
    .A( execution_unit_0.register_file_0.r1_5_ ),
    .B(_02566_),
    .C(_02636_),
    .Y(_02637_)
  );
  AOI22X1 _07903_ (
    .A( execution_unit_0.register_file_0.r10_5_ ),
    .B(_02583_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_5_ ),
    .Y(_02638_)
  );
  NAND2X1 _07904_ (
    .A(_02630_),
    .B(_02638_),
    .Y(_02639_)
  );
  AOI21X1 _07905_ (
    .A( execution_unit_0.register_file_0.r8_5_ ),
    .B(_02581_),
    .C(_02639_),
    .Y(_02640_)
  );
  OAI21X1 _07906_ (
    .A(_02560_),
    .B(_02592_),
    .C(_02633_),
    .Y(_02641_)
  );
  AOI22X1 _07907_ (
    .A( execution_unit_0.register_file_0.r6_5_ ),
    .B(_02575_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_5_ ),
    .Y(_02642_)
  );
  NAND2X1 _07908_ (
    .A(_02632_),
    .B(_02642_),
    .Y(_02643_)
  );
  NOR2X1 _07909_ (
    .A(_02641_),
    .B(_02643_),
    .Y(_02644_)
  );
  NAND2X1 _07910_ (
    .A(_02640_),
    .B(_02644_),
    .Y(_02645_)
  );
  NAND2X1 _07911_ (
    .A(_02631_),
    .B(_02637_),
    .Y(_02646_)
  );
  NOR2X1 _07912_ (
    .A(_02645_),
    .B(_02646_),
    .Y(_02647_)
  );
  INVX1 _07913_ (
    .A(_02647_),
    .Y( execution_unit_0.reg_src_5_ )
  );
  AOI22X1 _07914_ (
    .A( execution_unit_0.register_file_0.r10_6_ ),
    .B(_02583_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_6_ ),
    .Y(_02648_)
  );
  AOI22X1 _07915_ (
    .A( execution_unit_0.register_file_0.r3_6_ ),
    .B(_02574_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_6_ ),
    .Y(_02649_)
  );
  NAND2X1 _07916_ (
    .A(_02648_),
    .B(_02649_),
    .Y(_02650_)
  );
  AOI22X1 _07917_ (
    .A( execution_unit_0.register_file_0.r4_6_ ),
    .B(_02571_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_6_ ),
    .Y(_02651_)
  );
  AOI22X1 _07918_ (
    .A( execution_unit_0.register_file_0.r15_6_ ),
    .B(_02569_),
    .C(_02580_),
    .D( execution_unit_0.register_file_0.r14_6_ ),
    .Y(_02652_)
  );
  NAND2X1 _07919_ (
    .A(_02651_),
    .B(_02652_),
    .Y(_02653_)
  );
  NOR2X1 _07920_ (
    .A(_02650_),
    .B(_02653_),
    .Y(_02654_)
  );
  NAND2X1 _07921_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .B(_02572_),
    .Y(_02655_)
  );
  AOI22X1 _07922_ (
    .A( execution_unit_0.register_file_0.r1_6_ ),
    .B(_02566_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_6_ ),
    .Y(_02656_)
  );
  NAND2X1 _07923_ (
    .A(_02655_),
    .B(_02656_),
    .Y(_02657_)
  );
  AOI22X1 _07924_ (
    .A( execution_unit_0.register_file_0.r13_6_ ),
    .B(_02568_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_6_ ),
    .Y(_02658_)
  );
  AOI22X1 _07925_ (
    .A( execution_unit_0.register_file_0.r6_6_ ),
    .B(_02575_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_6_ ),
    .Y(_02659_)
  );
  NAND2X1 _07926_ (
    .A(_02658_),
    .B(_02659_),
    .Y(_02660_)
  );
  NOR2X1 _07927_ (
    .A(_02657_),
    .B(_02660_),
    .Y(_02661_)
  );
  NAND2X1 _07928_ (
    .A(_02654_),
    .B(_02661_),
    .Y( execution_unit_0.reg_src_6_ )
  );
  INVX1 _07929_ (
    .A( execution_unit_0.reg_src_6_ ),
    .Y(_02662_)
  );
  AOI22X1 _07930_ (
    .A( execution_unit_0.register_file_0.r15_7_ ),
    .B(_02569_),
    .C(_02571_),
    .D( execution_unit_0.register_file_0.r4_7_ ),
    .Y(_02663_)
  );
  AOI22X1 _07931_ (
    .A( execution_unit_0.register_file_0.r8_7_ ),
    .B(_02581_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_7_ ),
    .Y(_02664_)
  );
  NAND2X1 _07932_ (
    .A(_02663_),
    .B(_02664_),
    .Y(_02665_)
  );
  AOI22X1 _07933_ (
    .A( clock_module_0.scg1 ),
    .B(_02565_),
    .C(_02574_),
    .D( execution_unit_0.register_file_0.r3_7_ ),
    .Y(_02666_)
  );
  AOI22X1 _07934_ (
    .A( execution_unit_0.register_file_0.r13_7_ ),
    .B(_02568_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_7_ ),
    .Y(_02667_)
  );
  NAND2X1 _07935_ (
    .A(_02666_),
    .B(_02667_),
    .Y(_02668_)
  );
  NOR2X1 _07936_ (
    .A(_02665_),
    .B(_02668_),
    .Y(_02669_)
  );
  AOI22X1 _07937_ (
    .A( execution_unit_0.register_file_0.r6_7_ ),
    .B(_02575_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_7_ ),
    .Y(_02670_)
  );
  AOI22X1 _07938_ (
    .A( execution_unit_0.register_file_0.r1_7_ ),
    .B(_02566_),
    .C(_02572_),
    .D( dbg_0.UNUSED_pc_7_ ),
    .Y(_02671_)
  );
  NAND2X1 _07939_ (
    .A(_02670_),
    .B(_02671_),
    .Y(_02672_)
  );
  AOI22X1 _07940_ (
    .A( execution_unit_0.register_file_0.r5_7_ ),
    .B(_02589_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_7_ ),
    .Y(_02673_)
  );
  AOI22X1 _07941_ (
    .A( execution_unit_0.register_file_0.r14_7_ ),
    .B(_02580_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_7_ ),
    .Y(_02674_)
  );
  NAND2X1 _07942_ (
    .A(_02673_),
    .B(_02674_),
    .Y(_02675_)
  );
  NOR2X1 _07943_ (
    .A(_02672_),
    .B(_02675_),
    .Y(_02676_)
  );
  NAND2X1 _07944_ (
    .A(_02669_),
    .B(_02676_),
    .Y( execution_unit_0.reg_src_7_ )
  );
  INVX1 _07945_ (
    .A( execution_unit_0.reg_src_7_ ),
    .Y(_02677_)
  );
  NAND2X1 _07946_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_02678_)
  );
  INVX1 _07947_ (
    .A(_02678_),
    .Y( execution_unit_0.pc_sw_8_ )
  );
  AOI22X1 _07948_ (
    .A( execution_unit_0.register_file_0.r15_8_ ),
    .B(_02569_),
    .C(_02571_),
    .D( execution_unit_0.register_file_0.r4_8_ ),
    .Y(_02679_)
  );
  AOI22X1 _07949_ (
    .A( execution_unit_0.register_file_0.r8_8_ ),
    .B(_02581_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_8_ ),
    .Y(_02680_)
  );
  NAND2X1 _07950_ (
    .A(_02679_),
    .B(_02680_),
    .Y(_02681_)
  );
  AOI22X1 _07951_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .B(_02572_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_8_ ),
    .Y(_02682_)
  );
  AOI22X1 _07952_ (
    .A( execution_unit_0.register_file_0.r6_8_ ),
    .B(_02575_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_8_ ),
    .Y(_02683_)
  );
  NAND2X1 _07953_ (
    .A(_02682_),
    .B(_02683_),
    .Y(_02684_)
  );
  NOR2X1 _07954_ (
    .A(_02681_),
    .B(_02684_),
    .Y(_02685_)
  );
  AOI22X1 _07955_ (
    .A( execution_unit_0.register_file_0.r10_8_ ),
    .B(_02583_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_8_ ),
    .Y(_02686_)
  );
  AOI22X1 _07956_ (
    .A( execution_unit_0.alu_0.status_3_ ),
    .B(_02565_),
    .C(_02566_),
    .D( execution_unit_0.register_file_0.r1_8_ ),
    .Y(_02687_)
  );
  NAND2X1 _07957_ (
    .A(_02686_),
    .B(_02687_),
    .Y(_02688_)
  );
  AOI22X1 _07958_ (
    .A( execution_unit_0.register_file_0.r3_8_ ),
    .B(_02574_),
    .C(_02580_),
    .D( execution_unit_0.register_file_0.r14_8_ ),
    .Y(_02689_)
  );
  AOI22X1 _07959_ (
    .A( execution_unit_0.register_file_0.r13_8_ ),
    .B(_02568_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_8_ ),
    .Y(_02690_)
  );
  NAND2X1 _07960_ (
    .A(_02689_),
    .B(_02690_),
    .Y(_02691_)
  );
  NOR2X1 _07961_ (
    .A(_02688_),
    .B(_02691_),
    .Y(_02692_)
  );
  NAND2X1 _07962_ (
    .A(_02685_),
    .B(_02692_),
    .Y( execution_unit_0.reg_src_8_ )
  );
  INVX1 _07963_ (
    .A( execution_unit_0.reg_src_8_ ),
    .Y(_02693_)
  );
  AND2X1 _07964_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_9_ ),
    .Y( execution_unit_0.pc_sw_9_ )
  );
  INVX1 _07965_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .Y(_02694_)
  );
  NAND2X1 _07966_ (
    .A( execution_unit_0.register_file_0.r5_9_ ),
    .B(_02589_),
    .Y(_02695_)
  );
  NAND2X1 _07967_ (
    .A( execution_unit_0.register_file_0.r3_9_ ),
    .B(_02574_),
    .Y(_02696_)
  );
  AOI22X1 _07968_ (
    .A( execution_unit_0.register_file_0.r1_9_ ),
    .B(_02566_),
    .C(_02572_),
    .D( dbg_0.UNUSED_pc_9_ ),
    .Y(_02697_)
  );
  AOI22X1 _07969_ (
    .A( execution_unit_0.register_file_0.r15_9_ ),
    .B(_02569_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_9_ ),
    .Y(_02698_)
  );
  AOI22X1 _07970_ (
    .A( execution_unit_0.register_file_0.r14_9_ ),
    .B(_02580_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_9_ ),
    .Y(_02699_)
  );
  AOI22X1 _07971_ (
    .A( execution_unit_0.register_file_0.r6_9_ ),
    .B(_02575_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_9_ ),
    .Y(_02700_)
  );
  NAND2X1 _07972_ (
    .A(_02697_),
    .B(_02700_),
    .Y(_02701_)
  );
  AOI21X1 _07973_ (
    .A( execution_unit_0.register_file_0.r4_9_ ),
    .B(_02571_),
    .C(_02701_),
    .Y(_02702_)
  );
  AOI22X1 _07974_ (
    .A( execution_unit_0.register_file_0.r13_9_ ),
    .B(_02568_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_9_ ),
    .Y(_02703_)
  );
  NAND3X1 _07975_ (
    .A(_02695_),
    .B(_02696_),
    .C(_02703_),
    .Y(_02704_)
  );
  AOI22X1 _07976_ (
    .A( execution_unit_0.register_file_0.r9_9_ ),
    .B(_02588_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_9_ ),
    .Y(_02705_)
  );
  NAND3X1 _07977_ (
    .A(_02698_),
    .B(_02699_),
    .C(_02705_),
    .Y(_02706_)
  );
  NOR2X1 _07978_ (
    .A(_02704_),
    .B(_02706_),
    .Y(_02707_)
  );
  NAND2X1 _07979_ (
    .A(_02702_),
    .B(_02707_),
    .Y( execution_unit_0.reg_src_9_ )
  );
  INVX1 _07980_ (
    .A( execution_unit_0.reg_src_9_ ),
    .Y(_02708_)
  );
  NAND2X1 _07981_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_10_ ),
    .Y(_02709_)
  );
  INVX1 _07982_ (
    .A(_02709_),
    .Y( execution_unit_0.pc_sw_10_ )
  );
  AOI22X1 _07983_ (
    .A( execution_unit_0.register_file_0.r15_10_ ),
    .B(_02569_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_10_ ),
    .Y(_02710_)
  );
  AOI22X1 _07984_ (
    .A( dbg_0.UNUSED_pc_10_ ),
    .B(_02572_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_10_ ),
    .Y(_02711_)
  );
  NAND2X1 _07985_ (
    .A(_02710_),
    .B(_02711_),
    .Y(_02712_)
  );
  AOI22X1 _07986_ (
    .A( execution_unit_0.register_file_0.r1_10_ ),
    .B(_02566_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_10_ ),
    .Y(_02713_)
  );
  AOI22X1 _07987_ (
    .A( execution_unit_0.register_file_0.r13_10_ ),
    .B(_02568_),
    .C(_02580_),
    .D( execution_unit_0.register_file_0.r14_10_ ),
    .Y(_02714_)
  );
  NAND2X1 _07988_ (
    .A(_02713_),
    .B(_02714_),
    .Y(_02715_)
  );
  NOR2X1 _07989_ (
    .A(_02712_),
    .B(_02715_),
    .Y(_02716_)
  );
  NAND2X1 _07990_ (
    .A( execution_unit_0.register_file_0.r5_10_ ),
    .B(_02589_),
    .Y(_02717_)
  );
  AOI22X1 _07991_ (
    .A( execution_unit_0.register_file_0.r3_10_ ),
    .B(_02574_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_10_ ),
    .Y(_02718_)
  );
  NAND2X1 _07992_ (
    .A(_02717_),
    .B(_02718_),
    .Y(_02719_)
  );
  AOI22X1 _07993_ (
    .A( execution_unit_0.register_file_0.r4_10_ ),
    .B(_02571_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_10_ ),
    .Y(_02720_)
  );
  AOI22X1 _07994_ (
    .A( execution_unit_0.register_file_0.r6_10_ ),
    .B(_02575_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_10_ ),
    .Y(_02721_)
  );
  NAND2X1 _07995_ (
    .A(_02720_),
    .B(_02721_),
    .Y(_02722_)
  );
  NOR2X1 _07996_ (
    .A(_02719_),
    .B(_02722_),
    .Y(_02723_)
  );
  NAND2X1 _07997_ (
    .A(_02716_),
    .B(_02723_),
    .Y( execution_unit_0.reg_src_10_ )
  );
  INVX1 _07998_ (
    .A( execution_unit_0.reg_src_10_ ),
    .Y(_02724_)
  );
  AND2X1 _07999_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_11_ ),
    .Y( execution_unit_0.pc_sw_11_ )
  );
  INVX1 _08000_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .Y(_02725_)
  );
  NAND2X1 _08001_ (
    .A( execution_unit_0.register_file_0.r1_11_ ),
    .B(_02566_),
    .Y(_02726_)
  );
  AOI22X1 _08002_ (
    .A( execution_unit_0.register_file_0.r13_11_ ),
    .B(_02568_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_11_ ),
    .Y(_02727_)
  );
  AOI22X1 _08003_ (
    .A( execution_unit_0.register_file_0.r7_11_ ),
    .B(_02585_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_11_ ),
    .Y(_02728_)
  );
  AOI22X1 _08004_ (
    .A( execution_unit_0.register_file_0.r4_11_ ),
    .B(_02571_),
    .C(_02572_),
    .D( dbg_0.UNUSED_pc_11_ ),
    .Y(_02729_)
  );
  NAND2X1 _08005_ (
    .A(_02726_),
    .B(_02729_),
    .Y(_02730_)
  );
  AOI21X1 _08006_ (
    .A( execution_unit_0.register_file_0.r6_11_ ),
    .B(_02575_),
    .C(_02730_),
    .Y(_02731_)
  );
  AND2X1 _08007_ (
    .A(_02727_),
    .B(_02728_),
    .Y(_02732_)
  );
  AOI22X1 _08008_ (
    .A( execution_unit_0.register_file_0.r15_11_ ),
    .B(_02569_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_11_ ),
    .Y(_02733_)
  );
  AOI22X1 _08009_ (
    .A( execution_unit_0.register_file_0.r14_11_ ),
    .B(_02580_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_11_ ),
    .Y(_02734_)
  );
  AOI22X1 _08010_ (
    .A( execution_unit_0.register_file_0.r3_11_ ),
    .B(_02574_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_11_ ),
    .Y(_02735_)
  );
  NAND3X1 _08011_ (
    .A(_02733_),
    .B(_02734_),
    .C(_02735_),
    .Y(_02736_)
  );
  AOI21X1 _08012_ (
    .A( execution_unit_0.register_file_0.r11_11_ ),
    .B(_02591_),
    .C(_02736_),
    .Y(_02737_)
  );
  NAND3X1 _08013_ (
    .A(_02731_),
    .B(_02732_),
    .C(_02737_),
    .Y( execution_unit_0.reg_src_11_ )
  );
  INVX1 _08014_ (
    .A( execution_unit_0.reg_src_11_ ),
    .Y(_02738_)
  );
  NAND2X1 _08015_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_12_ ),
    .Y(_02739_)
  );
  INVX1 _08016_ (
    .A(_02739_),
    .Y( execution_unit_0.pc_sw_12_ )
  );
  AOI22X1 _08017_ (
    .A( execution_unit_0.register_file_0.r1_12_ ),
    .B(_02566_),
    .C(_02580_),
    .D( execution_unit_0.register_file_0.r14_12_ ),
    .Y(_02740_)
  );
  AOI22X1 _08018_ (
    .A( execution_unit_0.register_file_0.r3_12_ ),
    .B(_02574_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_12_ ),
    .Y(_02741_)
  );
  AND2X1 _08019_ (
    .A(_02740_),
    .B(_02741_),
    .Y(_02742_)
  );
  AOI22X1 _08020_ (
    .A( execution_unit_0.register_file_0.r11_12_ ),
    .B(_02591_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_12_ ),
    .Y(_02743_)
  );
  AOI22X1 _08021_ (
    .A( execution_unit_0.register_file_0.r7_12_ ),
    .B(_02585_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_12_ ),
    .Y(_02744_)
  );
  NAND3X1 _08022_ (
    .A(_02742_),
    .B(_02743_),
    .C(_02744_),
    .Y(_02745_)
  );
  AOI22X1 _08023_ (
    .A( execution_unit_0.register_file_0.r8_12_ ),
    .B(_02581_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_12_ ),
    .Y(_02746_)
  );
  INVX1 _08024_ (
    .A(_02746_),
    .Y(_02747_)
  );
  AOI21X1 _08025_ (
    .A( execution_unit_0.register_file_0.r4_12_ ),
    .B(_02571_),
    .C(_02747_),
    .Y(_02748_)
  );
  AOI22X1 _08026_ (
    .A( dbg_0.UNUSED_pc_12_ ),
    .B(_02572_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_12_ ),
    .Y(_02749_)
  );
  AOI22X1 _08027_ (
    .A( execution_unit_0.register_file_0.r13_12_ ),
    .B(_02568_),
    .C(_02569_),
    .D( execution_unit_0.register_file_0.r15_12_ ),
    .Y(_02750_)
  );
  NAND3X1 _08028_ (
    .A(_02748_),
    .B(_02749_),
    .C(_02750_),
    .Y(_02751_)
  );
  OR2X1 _08029_ (
    .A(_02745_),
    .B(_02751_),
    .Y( execution_unit_0.reg_src_12_ )
  );
  INVX1 _08030_ (
    .A( execution_unit_0.reg_src_12_ ),
    .Y(_02752_)
  );
  NAND2X1 _08031_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_13_ ),
    .Y(_02753_)
  );
  INVX1 _08032_ (
    .A(_02753_),
    .Y( execution_unit_0.pc_sw_13_ )
  );
  NAND2X1 _08033_ (
    .A( execution_unit_0.register_file_0.r4_13_ ),
    .B(_02571_),
    .Y(_02754_)
  );
  AOI22X1 _08034_ (
    .A( execution_unit_0.register_file_0.r1_13_ ),
    .B(_02566_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_13_ ),
    .Y(_02755_)
  );
  NAND2X1 _08035_ (
    .A(_02754_),
    .B(_02755_),
    .Y(_02756_)
  );
  AOI21X1 _08036_ (
    .A( execution_unit_0.register_file_0.r5_13_ ),
    .B(_02589_),
    .C(_02756_),
    .Y(_02757_)
  );
  AOI22X1 _08037_ (
    .A( dbg_0.UNUSED_pc_13_ ),
    .B(_02572_),
    .C(_02574_),
    .D( execution_unit_0.register_file_0.r3_13_ ),
    .Y(_02758_)
  );
  AOI22X1 _08038_ (
    .A( execution_unit_0.register_file_0.r8_13_ ),
    .B(_02581_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_13_ ),
    .Y(_02759_)
  );
  AND2X1 _08039_ (
    .A(_02758_),
    .B(_02759_),
    .Y(_02760_)
  );
  AOI22X1 _08040_ (
    .A( execution_unit_0.register_file_0.r15_13_ ),
    .B(_02569_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_13_ ),
    .Y(_02761_)
  );
  AOI22X1 _08041_ (
    .A( execution_unit_0.register_file_0.r13_13_ ),
    .B(_02568_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_13_ ),
    .Y(_02762_)
  );
  AOI22X1 _08042_ (
    .A( execution_unit_0.register_file_0.r14_13_ ),
    .B(_02580_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_13_ ),
    .Y(_02763_)
  );
  NAND3X1 _08043_ (
    .A(_02761_),
    .B(_02762_),
    .C(_02763_),
    .Y(_02764_)
  );
  AOI21X1 _08044_ (
    .A( execution_unit_0.register_file_0.r11_13_ ),
    .B(_02591_),
    .C(_02764_),
    .Y(_02765_)
  );
  NAND3X1 _08045_ (
    .A(_02757_),
    .B(_02760_),
    .C(_02765_),
    .Y( execution_unit_0.reg_src_13_ )
  );
  INVX1 _08046_ (
    .A( execution_unit_0.reg_src_13_ ),
    .Y(_02766_)
  );
  AND2X1 _08047_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_14_ ),
    .Y( execution_unit_0.pc_sw_14_ )
  );
  INVX1 _08048_ (
    .A( execution_unit_0.pc_sw_14_ ),
    .Y(_02767_)
  );
  NAND2X1 _08049_ (
    .A( execution_unit_0.register_file_0.r9_14_ ),
    .B(_02588_),
    .Y(_02768_)
  );
  AOI22X1 _08050_ (
    .A( execution_unit_0.register_file_0.r13_14_ ),
    .B(_02568_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_14_ ),
    .Y(_02769_)
  );
  AOI22X1 _08051_ (
    .A( execution_unit_0.register_file_0.r3_14_ ),
    .B(_02574_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_14_ ),
    .Y(_02770_)
  );
  AOI22X1 _08052_ (
    .A( execution_unit_0.register_file_0.r14_14_ ),
    .B(_02580_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_14_ ),
    .Y(_02771_)
  );
  NAND2X1 _08053_ (
    .A(_02769_),
    .B(_02771_),
    .Y(_02772_)
  );
  AOI21X1 _08054_ (
    .A( execution_unit_0.register_file_0.r10_14_ ),
    .B(_02583_),
    .C(_02772_),
    .Y(_02773_)
  );
  NAND2X1 _08055_ (
    .A(_02770_),
    .B(_02773_),
    .Y(_02774_)
  );
  AOI21X1 _08056_ (
    .A( execution_unit_0.register_file_0.r11_14_ ),
    .B(_02591_),
    .C(_02774_),
    .Y(_02775_)
  );
  AOI22X1 _08057_ (
    .A( execution_unit_0.register_file_0.r1_14_ ),
    .B(_02566_),
    .C(_02569_),
    .D( execution_unit_0.register_file_0.r15_14_ ),
    .Y(_02776_)
  );
  AOI22X1 _08058_ (
    .A( execution_unit_0.register_file_0.r8_14_ ),
    .B(_02581_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_14_ ),
    .Y(_02777_)
  );
  AOI22X1 _08059_ (
    .A( execution_unit_0.register_file_0.r4_14_ ),
    .B(_02571_),
    .C(_02572_),
    .D( dbg_0.UNUSED_pc_14_ ),
    .Y(_02778_)
  );
  NAND3X1 _08060_ (
    .A(_02768_),
    .B(_02777_),
    .C(_02778_),
    .Y(_02779_)
  );
  INVX1 _08061_ (
    .A(_02779_),
    .Y(_02780_)
  );
  NAND3X1 _08062_ (
    .A(_02775_),
    .B(_02776_),
    .C(_02780_),
    .Y( execution_unit_0.reg_src_14_ )
  );
  INVX1 _08063_ (
    .A( execution_unit_0.reg_src_14_ ),
    .Y(_02781_)
  );
  AND2X1 _08064_ (
    .A(_02544_),
    .B( execution_unit_0.alu_0.alu_out_15_ ),
    .Y( execution_unit_0.pc_sw_15_ )
  );
  INVX1 _08065_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .Y(_02782_)
  );
  AOI22X1 _08066_ (
    .A( execution_unit_0.register_file_0.r14_15_ ),
    .B(_02580_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_15_ ),
    .Y(_02783_)
  );
  AOI22X1 _08067_ (
    .A( execution_unit_0.register_file_0.r15_15_ ),
    .B(_02569_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_15_ ),
    .Y(_02784_)
  );
  AOI22X1 _08068_ (
    .A( execution_unit_0.register_file_0.r7_15_ ),
    .B(_02585_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_15_ ),
    .Y(_02785_)
  );
  OAI21X1 _08069_ (
    .A(_02564_),
    .B(_02576_),
    .C(_02785_),
    .Y(_02786_)
  );
  AOI21X1 _08070_ (
    .A( execution_unit_0.register_file_0.r9_15_ ),
    .B(_02588_),
    .C(_02786_),
    .Y(_02787_)
  );
  AND2X1 _08071_ (
    .A(_02783_),
    .B(_02784_),
    .Y(_02788_)
  );
  AOI22X1 _08072_ (
    .A( execution_unit_0.register_file_0.r13_15_ ),
    .B(_02568_),
    .C(_02574_),
    .D( execution_unit_0.register_file_0.r3_15_ ),
    .Y(_02789_)
  );
  AOI22X1 _08073_ (
    .A( dbg_0.UNUSED_pc_15_ ),
    .B(_02572_),
    .C(_02589_),
    .D( execution_unit_0.register_file_0.r5_15_ ),
    .Y(_02790_)
  );
  AOI22X1 _08074_ (
    .A( execution_unit_0.register_file_0.r4_15_ ),
    .B(_02571_),
    .C(_02581_),
    .D( execution_unit_0.register_file_0.r8_15_ ),
    .Y(_02791_)
  );
  NAND3X1 _08075_ (
    .A(_02789_),
    .B(_02790_),
    .C(_02791_),
    .Y(_02792_)
  );
  AOI21X1 _08076_ (
    .A( execution_unit_0.register_file_0.r1_15_ ),
    .B(_02566_),
    .C(_02792_),
    .Y(_02793_)
  );
  NAND3X1 _08077_ (
    .A(_02787_),
    .B(_02788_),
    .C(_02793_),
    .Y( execution_unit_0.reg_src_15_ )
  );
  INVX1 _08078_ (
    .A( execution_unit_0.reg_src_15_ ),
    .Y(_02794_)
  );
  AOI21X1 _08079_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_2_ ),
    .C( execution_unit_0.reg_sr_wr ),
    .Y(_02795_)
  );
  OAI21X1 _08080_ (
    .A(_02559_),
    .B(_02795_),
    .C(_02558_),
    .Y( clock_module_0.UNUSED_cpuoff )
  );
  MUX2X1 _08081_ (
    .A( execution_unit_0.register_file_0.r2_4_ ),
    .B( execution_unit_0.alu_0.alu_out_4_ ),
    .S(_02795_),
    .Y(_02796_)
  );
  NOR2X1 _08082_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B(_02796_),
    .Y(_01755_)
  );
  AOI21X1 _08083_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_0_ ),
    .C( execution_unit_0.reg_pc_call ),
    .Y(_02797_)
  );
  INVX1 _08084_ (
    .A(_02797_),
    .Y( execution_unit_0.pc_sw_wr )
  );
  NAND2X1 _08085_ (
    .A( execution_unit_0.register_file_0.r5_0_ ),
    .B(_02589_),
    .Y(_02798_)
  );
  AND2X1 _08086_ (
    .A( execution_unit_0.register_file_0.r8_0_ ),
    .B(_02581_),
    .Y(_02799_)
  );
  NAND3X1 _08087_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_4_ ),
    .C( execution_unit_0.register_file_0.r4_0_ ),
    .Y(_02800_)
  );
  NAND3X1 _08088_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_15_ ),
    .C( execution_unit_0.register_file_0.r15_0_ ),
    .Y(_02801_)
  );
  OAI21X1 _08089_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .C( execution_unit_0.alu_0.status_0_ ),
    .Y(_02802_)
  );
  NAND3X1 _08090_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_0_ ),
    .C( dbg_0.UNUSED_pc_0_ ),
    .Y(_02803_)
  );
  AND2X1 _08091_ (
    .A(_02802_),
    .B(_02803_),
    .Y(_02804_)
  );
  AOI22X1 _08092_ (
    .A( execution_unit_0.register_file_0.r13_0_ ),
    .B(_02568_),
    .C(_02583_),
    .D( execution_unit_0.register_file_0.r10_0_ ),
    .Y(_02805_)
  );
  NAND3X1 _08093_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_14_ ),
    .C( execution_unit_0.register_file_0.r14_0_ ),
    .Y(_02806_)
  );
  AOI22X1 _08094_ (
    .A( execution_unit_0.register_file_0.r3_0_ ),
    .B(_02574_),
    .C(_02575_),
    .D( execution_unit_0.register_file_0.r6_0_ ),
    .Y(_02807_)
  );
  NAND3X1 _08095_ (
    .A(_02798_),
    .B(_02804_),
    .C(_02807_),
    .Y(_02808_)
  );
  NAND3X1 _08096_ (
    .A(_02800_),
    .B(_02801_),
    .C(_02806_),
    .Y(_02809_)
  );
  OR2X1 _08097_ (
    .A(_02799_),
    .B(_02809_),
    .Y(_02810_)
  );
  AOI22X1 _08098_ (
    .A( execution_unit_0.register_file_0.r11_0_ ),
    .B(_02591_),
    .C(_02593_),
    .D( execution_unit_0.register_file_0.r12_0_ ),
    .Y(_02811_)
  );
  AOI22X1 _08099_ (
    .A( execution_unit_0.register_file_0.r7_0_ ),
    .B(_02585_),
    .C(_02588_),
    .D( execution_unit_0.register_file_0.r9_0_ ),
    .Y(_02812_)
  );
  NAND3X1 _08100_ (
    .A(_02805_),
    .B(_02811_),
    .C(_02812_),
    .Y(_02813_)
  );
  NOR3X1 _08101_ (
    .A(_02808_),
    .B(_02810_),
    .C(_02813_),
    .Y(_02814_)
  );
  INVX1 _08102_ (
    .A(_02814_),
    .Y( execution_unit_0.reg_src_0_ )
  );
  NAND3X1 _08103_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_14_ ),
    .C( execution_unit_0.register_file_0.r14_1_ ),
    .Y(_02815_)
  );
  NAND3X1 _08104_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_0_ ),
    .C( dbg_0.UNUSED_pc_1_ ),
    .Y(_02816_)
  );
  NAND2X1 _08105_ (
    .A(_02815_),
    .B(_02816_),
    .Y(_02817_)
  );
  NAND3X1 _08106_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_9_ ),
    .C( execution_unit_0.register_file_0.r9_1_ ),
    .Y(_02818_)
  );
  OAI21X1 _08107_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B( execution_unit_0.inst_src_2_ ),
    .C( execution_unit_0.alu_0.status_1_ ),
    .Y(_02819_)
  );
  NAND2X1 _08108_ (
    .A(_02818_),
    .B(_02819_),
    .Y(_02820_)
  );
  NOR2X1 _08109_ (
    .A(_02817_),
    .B(_02820_),
    .Y(_02821_)
  );
  NAND3X1 _08110_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_15_ ),
    .C( execution_unit_0.register_file_0.r15_1_ ),
    .Y(_02822_)
  );
  OAI21X1 _08111_ (
    .A(_02552_),
    .B(_02576_),
    .C(_02822_),
    .Y(_02823_)
  );
  NAND3X1 _08112_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_12_ ),
    .C( execution_unit_0.register_file_0.r12_1_ ),
    .Y(_02824_)
  );
  NAND3X1 _08113_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_1_ ),
    .C( execution_unit_0.register_file_0.r1_1_ ),
    .Y(_02825_)
  );
  NAND2X1 _08114_ (
    .A(_02824_),
    .B(_02825_),
    .Y(_02826_)
  );
  NOR2X1 _08115_ (
    .A(_02823_),
    .B(_02826_),
    .Y(_02827_)
  );
  AND2X1 _08116_ (
    .A(_02821_),
    .B(_02827_),
    .Y(_02828_)
  );
  NAND3X1 _08117_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_10_ ),
    .C( execution_unit_0.register_file_0.r10_1_ ),
    .Y(_02829_)
  );
  AOI22X1 _08118_ (
    .A( execution_unit_0.register_file_0.r10_1_ ),
    .B(_02583_),
    .C(_02591_),
    .D( execution_unit_0.register_file_0.r11_1_ ),
    .Y(_02830_)
  );
  NAND3X1 _08119_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_3_ ),
    .C( execution_unit_0.register_file_0.r3_1_ ),
    .Y(_02831_)
  );
  AOI22X1 _08120_ (
    .A( execution_unit_0.register_file_0.r3_1_ ),
    .B(_02574_),
    .C(_02585_),
    .D( execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02832_)
  );
  AND2X1 _08121_ (
    .A(_02830_),
    .B(_02832_),
    .Y(_02833_)
  );
  NAND3X1 _08122_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_8_ ),
    .C( execution_unit_0.register_file_0.r8_1_ ),
    .Y(_02834_)
  );
  NAND3X1 _08123_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_5_ ),
    .C( execution_unit_0.register_file_0.r5_1_ ),
    .Y(_02835_)
  );
  NAND2X1 _08124_ (
    .A(_02834_),
    .B(_02835_),
    .Y(_02836_)
  );
  NAND3X1 _08125_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_13_ ),
    .C( execution_unit_0.register_file_0.r13_1_ ),
    .Y(_02837_)
  );
  NAND3X1 _08126_ (
    .A(_02540_),
    .B( execution_unit_0.inst_src_4_ ),
    .C( execution_unit_0.register_file_0.r4_1_ ),
    .Y(_02838_)
  );
  NAND2X1 _08127_ (
    .A(_02837_),
    .B(_02838_),
    .Y(_02839_)
  );
  NOR2X1 _08128_ (
    .A(_02836_),
    .B(_02839_),
    .Y(_02840_)
  );
  AND2X1 _08129_ (
    .A(_02833_),
    .B(_02840_),
    .Y(_02841_)
  );
  NAND3X1 _08130_ (
    .A(_02818_),
    .B(_02819_),
    .C(_02831_),
    .Y(_02842_)
  );
  OAI21X1 _08131_ (
    .A(_02553_),
    .B(_02586_),
    .C(_02838_),
    .Y(_02843_)
  );
  NOR2X1 _08132_ (
    .A(_02842_),
    .B(_02843_),
    .Y(_02844_)
  );
  NAND3X1 _08133_ (
    .A(_02824_),
    .B(_02829_),
    .C(_02837_),
    .Y(_02845_)
  );
  AOI21X1 _08134_ (
    .A( execution_unit_0.register_file_0.r11_1_ ),
    .B(_02591_),
    .C(_02845_),
    .Y(_02846_)
  );
  NAND3X1 _08135_ (
    .A(_02816_),
    .B(_02825_),
    .C(_02835_),
    .Y(_02847_)
  );
  NAND2X1 _08136_ (
    .A(_02815_),
    .B(_02834_),
    .Y(_02848_)
  );
  NOR3X1 _08137_ (
    .A(_02823_),
    .B(_02847_),
    .C(_02848_),
    .Y(_02849_)
  );
  NAND3X1 _08138_ (
    .A(_02844_),
    .B(_02846_),
    .C(_02849_),
    .Y( execution_unit_0.reg_src_1_ )
  );
  AOI22X1 _08139_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_0_ ),
    .C( execution_unit_0.register_file_0.r14_0_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02850_)
  );
  NAND2X1 _08140_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_0_ ),
    .Y(_02851_)
  );
  AOI22X1 _08141_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_0_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_0_ ),
    .Y(_02852_)
  );
  AOI22X1 _08142_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.alu_0.status_0_ ),
    .C( execution_unit_0.register_file_0.r15_0_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02853_)
  );
  AND2X1 _08143_ (
    .A(_02852_),
    .B(_02853_),
    .Y(_02854_)
  );
  AOI22X1 _08144_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_0_ ),
    .C( execution_unit_0.register_file_0.r13_0_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02855_)
  );
  AOI22X1 _08145_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_0_ ),
    .C( execution_unit_0.register_file_0.r11_0_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02856_)
  );
  NAND3X1 _08146_ (
    .A(_02850_),
    .B(_02855_),
    .C(_02856_),
    .Y(_02857_)
  );
  AOI21X1 _08147_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_0_ ),
    .C(_02857_),
    .Y(_02858_)
  );
  AOI22X1 _08148_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_0_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_0_ ),
    .Y(_02859_)
  );
  NAND2X1 _08149_ (
    .A(_02851_),
    .B(_02859_),
    .Y(_02860_)
  );
  AOI21X1 _08150_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_0_ ),
    .C(_02860_),
    .Y(_02861_)
  );
  NAND3X1 _08151_ (
    .A(_02854_),
    .B(_02858_),
    .C(_02861_),
    .Y( dbg_0.dbg_reg_din_0_ )
  );
  AOI22X1 _08152_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_1_ ),
    .C( execution_unit_0.register_file_0.r4_1_ ),
    .D( execution_unit_0.inst_dest_4_ ),
    .Y(_02862_)
  );
  AOI22X1 _08153_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_1_ ),
    .C( execution_unit_0.register_file_0.r10_1_ ),
    .D( execution_unit_0.inst_dest_10_ ),
    .Y(_02863_)
  );
  NAND2X1 _08154_ (
    .A(_02862_),
    .B(_02863_),
    .Y(_02864_)
  );
  AOI22X1 _08155_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_1_ ),
    .C( execution_unit_0.register_file_0.r11_1_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02865_)
  );
  AOI22X1 _08156_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.alu_0.status_1_ ),
    .C( execution_unit_0.register_file_0.r14_1_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02866_)
  );
  NAND2X1 _08157_ (
    .A(_02865_),
    .B(_02866_),
    .Y(_02867_)
  );
  NOR2X1 _08158_ (
    .A(_02864_),
    .B(_02867_),
    .Y(_02868_)
  );
  AOI22X1 _08159_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_1_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_1_ ),
    .Y(_02869_)
  );
  AOI22X1 _08160_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_1_ ),
    .C( execution_unit_0.register_file_0.r15_1_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02870_)
  );
  NAND2X1 _08161_ (
    .A(_02869_),
    .B(_02870_),
    .Y(_02871_)
  );
  AOI22X1 _08162_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_1_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_1_ ),
    .Y(_02872_)
  );
  AOI22X1 _08163_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_1_ ),
    .C( execution_unit_0.register_file_0.r13_1_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02873_)
  );
  NAND2X1 _08164_ (
    .A(_02872_),
    .B(_02873_),
    .Y(_02874_)
  );
  NOR2X1 _08165_ (
    .A(_02871_),
    .B(_02874_),
    .Y(_02875_)
  );
  NAND2X1 _08166_ (
    .A(_02868_),
    .B(_02875_),
    .Y( dbg_0.dbg_reg_din_1_ )
  );
  AOI22X1 _08167_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_2_ ),
    .C( execution_unit_0.register_file_0.r8_2_ ),
    .D( execution_unit_0.inst_dest_8_ ),
    .Y(_02876_)
  );
  AOI22X1 _08168_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.alu_0.status_2_ ),
    .C( execution_unit_0.register_file_0.r14_2_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02877_)
  );
  NAND2X1 _08169_ (
    .A(_02876_),
    .B(_02877_),
    .Y(_02878_)
  );
  AOI22X1 _08170_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_2_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_2_ ),
    .Y(_02879_)
  );
  AOI22X1 _08171_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_2_ ),
    .C( execution_unit_0.register_file_0.r12_2_ ),
    .D( execution_unit_0.inst_dest_12_ ),
    .Y(_02880_)
  );
  NAND2X1 _08172_ (
    .A(_02879_),
    .B(_02880_),
    .Y(_02881_)
  );
  NOR2X1 _08173_ (
    .A(_02878_),
    .B(_02881_),
    .Y(_02882_)
  );
  AOI22X1 _08174_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_2_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_2_ ),
    .Y(_02883_)
  );
  AOI22X1 _08175_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_2_ ),
    .C( execution_unit_0.register_file_0.r15_2_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02884_)
  );
  NAND2X1 _08176_ (
    .A(_02883_),
    .B(_02884_),
    .Y(_02885_)
  );
  AOI22X1 _08177_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_2_ ),
    .C( execution_unit_0.register_file_0.r13_2_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02886_)
  );
  AOI22X1 _08178_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_2_ ),
    .C( execution_unit_0.register_file_0.r11_2_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02887_)
  );
  NAND2X1 _08179_ (
    .A(_02886_),
    .B(_02887_),
    .Y(_02888_)
  );
  NOR2X1 _08180_ (
    .A(_02885_),
    .B(_02888_),
    .Y(_02889_)
  );
  NAND2X1 _08181_ (
    .A(_02882_),
    .B(_02889_),
    .Y( dbg_0.dbg_reg_din_2_ )
  );
  AOI22X1 _08182_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_3_ ),
    .C( execution_unit_0.register_file_0.r7_3_ ),
    .D( execution_unit_0.inst_dest_7_ ),
    .Y(_02890_)
  );
  AOI22X1 _08183_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_3_ ),
    .C( execution_unit_0.register_file_0.r9_3_ ),
    .D( execution_unit_0.inst_dest_9_ ),
    .Y(_02891_)
  );
  NAND2X1 _08184_ (
    .A(_02890_),
    .B(_02891_),
    .Y(_02892_)
  );
  AOI22X1 _08185_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.gie ),
    .C( execution_unit_0.register_file_0.r3_3_ ),
    .D( execution_unit_0.inst_dest_3_ ),
    .Y(_02893_)
  );
  AOI22X1 _08186_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_3_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_3_ ),
    .Y(_02894_)
  );
  NAND2X1 _08187_ (
    .A(_02893_),
    .B(_02894_),
    .Y(_02895_)
  );
  NOR2X1 _08188_ (
    .A(_02892_),
    .B(_02895_),
    .Y(_02896_)
  );
  AOI22X1 _08189_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_3_ ),
    .C( execution_unit_0.register_file_0.r15_3_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02897_)
  );
  AOI22X1 _08190_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_3_ ),
    .C( execution_unit_0.register_file_0.r13_3_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02898_)
  );
  NAND2X1 _08191_ (
    .A(_02897_),
    .B(_02898_),
    .Y(_02899_)
  );
  AOI22X1 _08192_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_3_ ),
    .C( execution_unit_0.register_file_0.r14_3_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02900_)
  );
  AOI22X1 _08193_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_3_ ),
    .C( execution_unit_0.register_file_0.r11_3_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02901_)
  );
  NAND2X1 _08194_ (
    .A(_02900_),
    .B(_02901_),
    .Y(_02902_)
  );
  NOR2X1 _08195_ (
    .A(_02899_),
    .B(_02902_),
    .Y(_02903_)
  );
  NAND2X1 _08196_ (
    .A(_02896_),
    .B(_02903_),
    .Y( dbg_0.dbg_reg_din_3_ )
  );
  AOI22X1 _08197_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_4_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_4_ ),
    .Y(_02904_)
  );
  AOI22X1 _08198_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_4_ ),
    .C( execution_unit_0.register_file_0.r8_4_ ),
    .D( execution_unit_0.inst_dest_8_ ),
    .Y(_02905_)
  );
  NAND2X1 _08199_ (
    .A(_02904_),
    .B(_02905_),
    .Y(_01987_)
  );
  AOI22X1 _08200_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_4_ ),
    .C( execution_unit_0.register_file_0.r12_4_ ),
    .D( execution_unit_0.inst_dest_12_ ),
    .Y(_01988_)
  );
  AOI22X1 _08201_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_4_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_4_ ),
    .Y(_01989_)
  );
  NAND2X1 _08202_ (
    .A(_01988_),
    .B(_01989_),
    .Y(_01990_)
  );
  NOR2X1 _08203_ (
    .A(_01987_),
    .B(_01990_),
    .Y(_01991_)
  );
  AOI22X1 _08204_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_4_ ),
    .C( execution_unit_0.register_file_0.r13_4_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_01992_)
  );
  AOI22X1 _08205_ (
    .A( execution_unit_0.inst_dest_11_ ),
    .B( execution_unit_0.register_file_0.r11_4_ ),
    .C( execution_unit_0.register_file_0.r15_4_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_01993_)
  );
  NAND2X1 _08206_ (
    .A(_01992_),
    .B(_01993_),
    .Y(_01994_)
  );
  AOI22X1 _08207_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.register_file_0.r2_4_ ),
    .C( execution_unit_0.register_file_0.r6_4_ ),
    .D( execution_unit_0.inst_dest_6_ ),
    .Y(_01995_)
  );
  AOI22X1 _08208_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_4_ ),
    .C( execution_unit_0.register_file_0.r14_4_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_01996_)
  );
  NAND2X1 _08209_ (
    .A(_01995_),
    .B(_01996_),
    .Y(_01997_)
  );
  NOR2X1 _08210_ (
    .A(_01994_),
    .B(_01997_),
    .Y(_01998_)
  );
  NAND2X1 _08211_ (
    .A(_01991_),
    .B(_01998_),
    .Y( dbg_0.dbg_reg_din_4_ )
  );
  AOI22X1 _08212_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( clock_module_0.oscoff ),
    .C( execution_unit_0.register_file_0.r13_5_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_01999_)
  );
  AOI22X1 _08213_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_5_ ),
    .C( execution_unit_0.register_file_0.r10_5_ ),
    .D( execution_unit_0.inst_dest_10_ ),
    .Y(_02000_)
  );
  NAND2X1 _08214_ (
    .A(_01999_),
    .B(_02000_),
    .Y(_02001_)
  );
  AOI22X1 _08215_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_5_ ),
    .C( execution_unit_0.register_file_0.r9_5_ ),
    .D( execution_unit_0.inst_dest_9_ ),
    .Y(_02002_)
  );
  AOI22X1 _08216_ (
    .A( execution_unit_0.inst_dest_11_ ),
    .B( execution_unit_0.register_file_0.r11_5_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_5_ ),
    .Y(_02003_)
  );
  NAND2X1 _08217_ (
    .A(_02002_),
    .B(_02003_),
    .Y(_02004_)
  );
  NOR2X1 _08218_ (
    .A(_02001_),
    .B(_02004_),
    .Y(_02005_)
  );
  AOI22X1 _08219_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_5_ ),
    .C( execution_unit_0.register_file_0.r14_5_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02006_)
  );
  AOI22X1 _08220_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_5_ ),
    .C( execution_unit_0.register_file_0.r6_5_ ),
    .D( execution_unit_0.inst_dest_6_ ),
    .Y(_02007_)
  );
  NAND2X1 _08221_ (
    .A(_02006_),
    .B(_02007_),
    .Y(_02008_)
  );
  AOI22X1 _08222_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_5_ ),
    .C( execution_unit_0.register_file_0.r8_5_ ),
    .D( execution_unit_0.inst_dest_8_ ),
    .Y(_02009_)
  );
  AOI22X1 _08223_ (
    .A( execution_unit_0.inst_dest_15_ ),
    .B( execution_unit_0.register_file_0.r15_5_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_5_ ),
    .Y(_02010_)
  );
  NAND2X1 _08224_ (
    .A(_02009_),
    .B(_02010_),
    .Y(_02011_)
  );
  NOR2X1 _08225_ (
    .A(_02008_),
    .B(_02011_),
    .Y(_02012_)
  );
  NAND2X1 _08226_ (
    .A(_02005_),
    .B(_02012_),
    .Y( dbg_0.dbg_reg_din_5_ )
  );
  AOI22X1 _08227_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_6_ ),
    .C( execution_unit_0.register_file_0.r9_6_ ),
    .D( execution_unit_0.inst_dest_9_ ),
    .Y(_02013_)
  );
  AOI22X1 _08228_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_6_ ),
    .C( execution_unit_0.register_file_0.r14_6_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02014_)
  );
  NAND2X1 _08229_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_6_ ),
    .Y(_02015_)
  );
  NAND2X1 _08230_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .B( execution_unit_0.inst_dest_0_ ),
    .Y(_02016_)
  );
  AOI22X1 _08231_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_6_ ),
    .C( execution_unit_0.register_file_0.r5_6_ ),
    .D( execution_unit_0.inst_dest_5_ ),
    .Y(_02017_)
  );
  AOI22X1 _08232_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_6_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_6_ ),
    .Y(_02018_)
  );
  NAND2X1 _08233_ (
    .A(_02017_),
    .B(_02018_),
    .Y(_02019_)
  );
  AOI21X1 _08234_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_6_ ),
    .C(_02019_),
    .Y(_02020_)
  );
  NAND3X1 _08235_ (
    .A(_02014_),
    .B(_02015_),
    .C(_02016_),
    .Y(_02021_)
  );
  AOI22X1 _08236_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_6_ ),
    .C( execution_unit_0.register_file_0.r15_6_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02022_)
  );
  AOI22X1 _08237_ (
    .A( execution_unit_0.inst_dest_11_ ),
    .B( execution_unit_0.register_file_0.r11_6_ ),
    .C( execution_unit_0.register_file_0.r13_6_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02023_)
  );
  NAND3X1 _08238_ (
    .A(_02013_),
    .B(_02022_),
    .C(_02023_),
    .Y(_02024_)
  );
  NOR2X1 _08239_ (
    .A(_02021_),
    .B(_02024_),
    .Y(_02025_)
  );
  NAND2X1 _08240_ (
    .A(_02020_),
    .B(_02025_),
    .Y( dbg_0.dbg_reg_din_6_ )
  );
  AOI22X1 _08241_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_7_ ),
    .C( execution_unit_0.register_file_0.r12_7_ ),
    .D( execution_unit_0.inst_dest_12_ ),
    .Y(_02026_)
  );
  AOI22X1 _08242_ (
    .A( execution_unit_0.inst_dest_11_ ),
    .B( execution_unit_0.register_file_0.r11_7_ ),
    .C( execution_unit_0.register_file_0.r13_7_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02027_)
  );
  NAND2X1 _08243_ (
    .A(_02026_),
    .B(_02027_),
    .Y(_02028_)
  );
  AOI22X1 _08244_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_7_ ),
    .C( execution_unit_0.register_file_0.r14_7_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02029_)
  );
  AOI22X1 _08245_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_7_ ),
    .C( execution_unit_0.register_file_0.r5_7_ ),
    .D( execution_unit_0.inst_dest_5_ ),
    .Y(_02030_)
  );
  NAND2X1 _08246_ (
    .A(_02029_),
    .B(_02030_),
    .Y(_02031_)
  );
  NOR2X1 _08247_ (
    .A(_02028_),
    .B(_02031_),
    .Y(_02032_)
  );
  AOI22X1 _08248_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_7_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_7_ ),
    .Y(_02033_)
  );
  AOI22X1 _08249_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( clock_module_0.scg1 ),
    .C( execution_unit_0.register_file_0.r15_7_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02034_)
  );
  NAND2X1 _08250_ (
    .A(_02033_),
    .B(_02034_),
    .Y(_02035_)
  );
  AOI22X1 _08251_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_7_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_7_ ),
    .Y(_02036_)
  );
  AOI22X1 _08252_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_7_ ),
    .C( execution_unit_0.register_file_0.r10_7_ ),
    .D( execution_unit_0.inst_dest_10_ ),
    .Y(_02037_)
  );
  NAND2X1 _08253_ (
    .A(_02036_),
    .B(_02037_),
    .Y(_02038_)
  );
  NOR2X1 _08254_ (
    .A(_02035_),
    .B(_02038_),
    .Y(_02039_)
  );
  NAND2X1 _08255_ (
    .A(_02032_),
    .B(_02039_),
    .Y( dbg_0.dbg_reg_din_7_ )
  );
  AOI22X1 _08256_ (
    .A( execution_unit_0.inst_dest_2_ ),
    .B( execution_unit_0.alu_0.status_3_ ),
    .C( execution_unit_0.register_file_0.r10_8_ ),
    .D( execution_unit_0.inst_dest_10_ ),
    .Y(_02040_)
  );
  AOI22X1 _08257_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_8_ ),
    .C( execution_unit_0.register_file_0.r13_8_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02041_)
  );
  NAND2X1 _08258_ (
    .A(_02040_),
    .B(_02041_),
    .Y(_02042_)
  );
  AOI22X1 _08259_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_8_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_8_ ),
    .Y(_02043_)
  );
  AOI22X1 _08260_ (
    .A( execution_unit_0.inst_dest_14_ ),
    .B( execution_unit_0.register_file_0.r14_8_ ),
    .C( execution_unit_0.register_file_0.r15_8_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02044_)
  );
  NAND2X1 _08261_ (
    .A(_02043_),
    .B(_02044_),
    .Y(_02045_)
  );
  NOR2X1 _08262_ (
    .A(_02042_),
    .B(_02045_),
    .Y(_02046_)
  );
  AOI22X1 _08263_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_8_ ),
    .C( execution_unit_0.register_file_0.r12_8_ ),
    .D( execution_unit_0.inst_dest_12_ ),
    .Y(_02047_)
  );
  AOI22X1 _08264_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_8_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_8_ ),
    .Y(_02048_)
  );
  NAND2X1 _08265_ (
    .A(_02047_),
    .B(_02048_),
    .Y(_02049_)
  );
  AOI22X1 _08266_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_8_ ),
    .C( execution_unit_0.register_file_0.r11_8_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02050_)
  );
  AOI22X1 _08267_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_8_ ),
    .C( execution_unit_0.register_file_0.r8_8_ ),
    .D( execution_unit_0.inst_dest_8_ ),
    .Y(_02051_)
  );
  NAND2X1 _08268_ (
    .A(_02050_),
    .B(_02051_),
    .Y(_02052_)
  );
  NOR2X1 _08269_ (
    .A(_02049_),
    .B(_02052_),
    .Y(_02053_)
  );
  NAND2X1 _08270_ (
    .A(_02046_),
    .B(_02053_),
    .Y( dbg_0.dbg_reg_din_8_ )
  );
  NAND2X1 _08271_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_9_ ),
    .Y(_02054_)
  );
  NAND2X1 _08272_ (
    .A( execution_unit_0.inst_dest_15_ ),
    .B( execution_unit_0.register_file_0.r15_9_ ),
    .Y(_02055_)
  );
  AOI22X1 _08273_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_9_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_9_ ),
    .Y(_02056_)
  );
  AOI22X1 _08274_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_9_ ),
    .C( execution_unit_0.register_file_0.r8_9_ ),
    .D( execution_unit_0.inst_dest_8_ ),
    .Y(_02057_)
  );
  NAND2X1 _08275_ (
    .A(_02054_),
    .B(_02057_),
    .Y(_02058_)
  );
  AOI22X1 _08276_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_9_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_9_ ),
    .Y(_02059_)
  );
  NAND2X1 _08277_ (
    .A(_02055_),
    .B(_02059_),
    .Y(_02060_)
  );
  NOR2X1 _08278_ (
    .A(_02058_),
    .B(_02060_),
    .Y(_02061_)
  );
  AOI22X1 _08279_ (
    .A( execution_unit_0.inst_dest_13_ ),
    .B( execution_unit_0.register_file_0.r13_9_ ),
    .C( execution_unit_0.register_file_0.r14_9_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02062_)
  );
  AOI22X1 _08280_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_9_ ),
    .C( execution_unit_0.register_file_0.r12_9_ ),
    .D( execution_unit_0.inst_dest_12_ ),
    .Y(_02063_)
  );
  AOI22X1 _08281_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_9_ ),
    .C( execution_unit_0.register_file_0.r11_9_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02064_)
  );
  NAND3X1 _08282_ (
    .A(_02062_),
    .B(_02063_),
    .C(_02064_),
    .Y(_02065_)
  );
  AOI21X1 _08283_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_9_ ),
    .C(_02065_),
    .Y(_02066_)
  );
  NAND3X1 _08284_ (
    .A(_02056_),
    .B(_02061_),
    .C(_02066_),
    .Y( dbg_0.dbg_reg_din_9_ )
  );
  AOI22X1 _08285_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_10_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_10_ ),
    .Y(_02067_)
  );
  AOI22X1 _08286_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_10_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_10_ ),
    .Y(_02068_)
  );
  AND2X1 _08287_ (
    .A(_02067_),
    .B(_02068_),
    .Y(_02069_)
  );
  AOI22X1 _08288_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_10_ ),
    .C( execution_unit_0.register_file_0.r14_10_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02070_)
  );
  AOI22X1 _08289_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_10_ ),
    .C( execution_unit_0.register_file_0.r15_10_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02071_)
  );
  NAND3X1 _08290_ (
    .A(_02069_),
    .B(_02070_),
    .C(_02071_),
    .Y(_02072_)
  );
  AOI22X1 _08291_ (
    .A( execution_unit_0.inst_dest_11_ ),
    .B( execution_unit_0.register_file_0.r11_10_ ),
    .C( execution_unit_0.register_file_0.r13_10_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02073_)
  );
  INVX1 _08292_ (
    .A(_02073_),
    .Y(_02074_)
  );
  AOI21X1 _08293_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_10_ ),
    .C(_02074_),
    .Y(_02075_)
  );
  AOI22X1 _08294_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_10_ ),
    .C( execution_unit_0.register_file_0.r9_10_ ),
    .D( execution_unit_0.inst_dest_9_ ),
    .Y(_02076_)
  );
  AOI22X1 _08295_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_10_ ),
    .C( execution_unit_0.register_file_0.r6_10_ ),
    .D( execution_unit_0.inst_dest_6_ ),
    .Y(_02077_)
  );
  NAND3X1 _08296_ (
    .A(_02075_),
    .B(_02076_),
    .C(_02077_),
    .Y(_02078_)
  );
  OR2X1 _08297_ (
    .A(_02072_),
    .B(_02078_),
    .Y( dbg_0.dbg_reg_din_10_ )
  );
  NAND2X1 _08298_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_11_ ),
    .Y(_02079_)
  );
  NAND2X1 _08299_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_11_ ),
    .Y(_02080_)
  );
  AOI22X1 _08300_ (
    .A( execution_unit_0.inst_dest_13_ ),
    .B( execution_unit_0.register_file_0.r13_11_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_11_ ),
    .Y(_02081_)
  );
  NAND2X1 _08301_ (
    .A(_02079_),
    .B(_02081_),
    .Y(_02082_)
  );
  AOI21X1 _08302_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_11_ ),
    .C(_02082_),
    .Y(_02083_)
  );
  AOI22X1 _08303_ (
    .A( execution_unit_0.inst_dest_14_ ),
    .B( execution_unit_0.register_file_0.r14_11_ ),
    .C( execution_unit_0.register_file_0.r15_11_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02084_)
  );
  AOI22X1 _08304_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_11_ ),
    .C( execution_unit_0.register_file_0.r11_11_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02085_)
  );
  NAND2X1 _08305_ (
    .A(_02084_),
    .B(_02085_),
    .Y(_02086_)
  );
  AOI21X1 _08306_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_11_ ),
    .C(_02086_),
    .Y(_02087_)
  );
  AOI22X1 _08307_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_11_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_11_ ),
    .Y(_02088_)
  );
  AOI22X1 _08308_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_11_ ),
    .C( execution_unit_0.register_file_0.r8_11_ ),
    .D( execution_unit_0.inst_dest_8_ ),
    .Y(_02089_)
  );
  NAND3X1 _08309_ (
    .A(_02080_),
    .B(_02088_),
    .C(_02089_),
    .Y(_02090_)
  );
  AOI21X1 _08310_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_11_ ),
    .C(_02090_),
    .Y(_02091_)
  );
  NAND3X1 _08311_ (
    .A(_02083_),
    .B(_02087_),
    .C(_02091_),
    .Y( dbg_0.dbg_reg_din_11_ )
  );
  NAND2X1 _08312_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_12_ ),
    .Y(_02092_)
  );
  NAND2X1 _08313_ (
    .A( dbg_0.UNUSED_pc_12_ ),
    .B( execution_unit_0.inst_dest_0_ ),
    .Y(_02093_)
  );
  AOI22X1 _08314_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_12_ ),
    .C( execution_unit_0.register_file_0.r14_12_ ),
    .D( execution_unit_0.inst_dest_14_ ),
    .Y(_02094_)
  );
  NAND2X1 _08315_ (
    .A(_02093_),
    .B(_02094_),
    .Y(_02095_)
  );
  AOI21X1 _08316_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_12_ ),
    .C(_02095_),
    .Y(_02096_)
  );
  AOI22X1 _08317_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_12_ ),
    .C( execution_unit_0.register_file_0.r5_12_ ),
    .D( execution_unit_0.inst_dest_5_ ),
    .Y(_02097_)
  );
  AOI22X1 _08318_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_12_ ),
    .C( execution_unit_0.register_file_0.r3_12_ ),
    .D( execution_unit_0.inst_dest_3_ ),
    .Y(_02098_)
  );
  NAND2X1 _08319_ (
    .A(_02097_),
    .B(_02098_),
    .Y(_02099_)
  );
  AOI21X1 _08320_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_12_ ),
    .C(_02099_),
    .Y(_02100_)
  );
  AOI22X1 _08321_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_12_ ),
    .C( execution_unit_0.register_file_0.r15_12_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02101_)
  );
  AOI22X1 _08322_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_12_ ),
    .C( execution_unit_0.register_file_0.r11_12_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02102_)
  );
  NAND3X1 _08323_ (
    .A(_02092_),
    .B(_02101_),
    .C(_02102_),
    .Y(_02103_)
  );
  AOI21X1 _08324_ (
    .A( execution_unit_0.inst_dest_13_ ),
    .B( execution_unit_0.register_file_0.r13_12_ ),
    .C(_02103_),
    .Y(_02104_)
  );
  NAND3X1 _08325_ (
    .A(_02096_),
    .B(_02100_),
    .C(_02104_),
    .Y( dbg_0.dbg_reg_din_12_ )
  );
  AOI22X1 _08326_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_13_ ),
    .C( execution_unit_0.register_file_0.r11_13_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02105_)
  );
  AOI22X1 _08327_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_13_ ),
    .C( execution_unit_0.register_file_0.r5_13_ ),
    .D( execution_unit_0.inst_dest_5_ ),
    .Y(_02106_)
  );
  AND2X1 _08328_ (
    .A(_02105_),
    .B(_02106_),
    .Y(_02107_)
  );
  AOI22X1 _08329_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_13_ ),
    .C( execution_unit_0.register_file_0.r13_13_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02108_)
  );
  AOI22X1 _08330_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_13_ ),
    .C( execution_unit_0.register_file_0.r9_13_ ),
    .D( execution_unit_0.inst_dest_9_ ),
    .Y(_02109_)
  );
  NAND3X1 _08331_ (
    .A(_02107_),
    .B(_02108_),
    .C(_02109_),
    .Y(_02110_)
  );
  AOI22X1 _08332_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_13_ ),
    .C( execution_unit_0.register_file_0.r10_13_ ),
    .D( execution_unit_0.inst_dest_10_ ),
    .Y(_02111_)
  );
  INVX1 _08333_ (
    .A(_02111_),
    .Y(_02112_)
  );
  AOI21X1 _08334_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_13_ ),
    .C(_02112_),
    .Y(_02113_)
  );
  AOI22X1 _08335_ (
    .A( execution_unit_0.inst_dest_14_ ),
    .B( execution_unit_0.register_file_0.r14_13_ ),
    .C( execution_unit_0.register_file_0.r15_13_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02114_)
  );
  AOI22X1 _08336_ (
    .A( dbg_0.UNUSED_pc_13_ ),
    .B( execution_unit_0.inst_dest_0_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_13_ ),
    .Y(_02115_)
  );
  NAND3X1 _08337_ (
    .A(_02113_),
    .B(_02114_),
    .C(_02115_),
    .Y(_02116_)
  );
  OR2X1 _08338_ (
    .A(_02110_),
    .B(_02116_),
    .Y( dbg_0.dbg_reg_din_13_ )
  );
  AOI22X1 _08339_ (
    .A( execution_unit_0.inst_dest_9_ ),
    .B( execution_unit_0.register_file_0.r9_14_ ),
    .C( execution_unit_0.register_file_0.r15_14_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02117_)
  );
  NAND2X1 _08340_ (
    .A( execution_unit_0.inst_dest_12_ ),
    .B( execution_unit_0.register_file_0.r12_14_ ),
    .Y(_02118_)
  );
  NAND2X1 _08341_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_14_ ),
    .Y(_02119_)
  );
  AOI22X1 _08342_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_14_ ),
    .C( execution_unit_0.register_file_0.r13_14_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02120_)
  );
  NAND2X1 _08343_ (
    .A(_02118_),
    .B(_02120_),
    .Y(_02121_)
  );
  AOI22X1 _08344_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_14_ ),
    .C( execution_unit_0.register_file_0.r6_14_ ),
    .D( execution_unit_0.inst_dest_6_ ),
    .Y(_02122_)
  );
  AOI22X1 _08345_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_14_ ),
    .C( execution_unit_0.register_file_0.r5_14_ ),
    .D( execution_unit_0.inst_dest_5_ ),
    .Y(_02123_)
  );
  AOI22X1 _08346_ (
    .A( dbg_0.UNUSED_pc_14_ ),
    .B( execution_unit_0.inst_dest_0_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_14_ ),
    .Y(_02124_)
  );
  NAND3X1 _08347_ (
    .A(_02122_),
    .B(_02123_),
    .C(_02124_),
    .Y(_02125_)
  );
  AOI21X1 _08348_ (
    .A( execution_unit_0.inst_dest_14_ ),
    .B( execution_unit_0.register_file_0.r14_14_ ),
    .C(_02125_),
    .Y(_02126_)
  );
  AOI22X1 _08349_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_14_ ),
    .C( execution_unit_0.register_file_0.r11_14_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02127_)
  );
  NAND2X1 _08350_ (
    .A(_02119_),
    .B(_02127_),
    .Y(_02128_)
  );
  NOR2X1 _08351_ (
    .A(_02121_),
    .B(_02128_),
    .Y(_02129_)
  );
  NAND3X1 _08352_ (
    .A(_02117_),
    .B(_02126_),
    .C(_02129_),
    .Y( dbg_0.dbg_reg_din_14_ )
  );
  AOI22X1 _08353_ (
    .A( execution_unit_0.inst_dest_14_ ),
    .B( execution_unit_0.register_file_0.r14_15_ ),
    .C( execution_unit_0.inst_dest_3_ ),
    .D( execution_unit_0.register_file_0.r3_15_ ),
    .Y(_02130_)
  );
  AOI22X1 _08354_ (
    .A( execution_unit_0.inst_dest_8_ ),
    .B( execution_unit_0.register_file_0.r8_15_ ),
    .C( execution_unit_0.register_file_0.r15_15_ ),
    .D( execution_unit_0.inst_dest_15_ ),
    .Y(_02131_)
  );
  AND2X1 _08355_ (
    .A(_02130_),
    .B(_02131_),
    .Y(_02132_)
  );
  AOI22X1 _08356_ (
    .A( execution_unit_0.inst_dest_10_ ),
    .B( execution_unit_0.register_file_0.r10_15_ ),
    .C( execution_unit_0.register_file_0.r13_15_ ),
    .D( execution_unit_0.inst_dest_13_ ),
    .Y(_02133_)
  );
  AOI22X1 _08357_ (
    .A( execution_unit_0.inst_dest_7_ ),
    .B( execution_unit_0.register_file_0.r7_15_ ),
    .C( execution_unit_0.register_file_0.r9_15_ ),
    .D( execution_unit_0.inst_dest_9_ ),
    .Y(_02134_)
  );
  NAND3X1 _08358_ (
    .A(_02132_),
    .B(_02133_),
    .C(_02134_),
    .Y(_02135_)
  );
  AOI22X1 _08359_ (
    .A( execution_unit_0.inst_dest_5_ ),
    .B( execution_unit_0.register_file_0.r5_15_ ),
    .C( execution_unit_0.register_file_0.r12_15_ ),
    .D( execution_unit_0.inst_dest_12_ ),
    .Y(_02136_)
  );
  INVX1 _08360_ (
    .A(_02136_),
    .Y(_02137_)
  );
  AOI21X1 _08361_ (
    .A( execution_unit_0.inst_dest_4_ ),
    .B( execution_unit_0.register_file_0.r4_15_ ),
    .C(_02137_),
    .Y(_02138_)
  );
  AOI22X1 _08362_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.register_file_0.r1_15_ ),
    .C( execution_unit_0.register_file_0.r11_15_ ),
    .D( execution_unit_0.inst_dest_11_ ),
    .Y(_02139_)
  );
  AOI22X1 _08363_ (
    .A( execution_unit_0.inst_dest_6_ ),
    .B( execution_unit_0.register_file_0.r6_15_ ),
    .C( execution_unit_0.inst_dest_0_ ),
    .D( dbg_0.UNUSED_pc_15_ ),
    .Y(_02140_)
  );
  NAND3X1 _08364_ (
    .A(_02138_),
    .B(_02139_),
    .C(_02140_),
    .Y(_02141_)
  );
  OR2X1 _08365_ (
    .A(_02135_),
    .B(_02141_),
    .Y( dbg_0.dbg_reg_din_15_ )
  );
  MUX2X1 _08366_ (
    .A( execution_unit_0.alu_0.status_1_ ),
    .B( execution_unit_0.alu_0.alu_out_1_ ),
    .S(_02795_),
    .Y(_02142_)
  );
  OAI21X1 _08367_ (
    .A(_02542_),
    .B( execution_unit_0.alu_0.Z ),
    .C(_02540_),
    .Y(_02143_)
  );
  AOI21X1 _08368_ (
    .A(_02542_),
    .B(_02142_),
    .C(_02143_),
    .Y(_01757_)
  );
  MUX2X1 _08369_ (
    .A( execution_unit_0.alu_0.status_2_ ),
    .B( execution_unit_0.alu_0.alu_out_2_ ),
    .S(_02795_),
    .Y(_02144_)
  );
  OAI21X1 _08370_ (
    .A(_02543_),
    .B( execution_unit_0.alu_0.N ),
    .C(_02540_),
    .Y(_02145_)
  );
  AOI21X1 _08371_ (
    .A(_02543_),
    .B(_02144_),
    .C(_02145_),
    .Y(_01758_)
  );
  AND2X1 _08372_ (
    .A(_02540_),
    .B(_02795_),
    .Y(_02146_)
  );
  NAND2X1 _08373_ (
    .A( execution_unit_0.gie ),
    .B(_02146_),
    .Y(_02147_)
  );
  NAND2X1 _08374_ (
    .A(_02540_),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_02148_)
  );
  OAI21X1 _08375_ (
    .A(_02795_),
    .B(_02148_),
    .C(_02147_),
    .Y(_01759_)
  );
  NAND2X1 _08376_ (
    .A( clock_module_0.oscoff ),
    .B(_02146_),
    .Y(_02149_)
  );
  NAND2X1 _08377_ (
    .A(_02540_),
    .B( execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_02150_)
  );
  OAI21X1 _08378_ (
    .A(_02795_),
    .B(_02150_),
    .C(_02149_),
    .Y(_01760_)
  );
  NAND2X1 _08379_ (
    .A( clock_module_0.scg1 ),
    .B(_02146_),
    .Y(_02151_)
  );
  NAND2X1 _08380_ (
    .A(_02540_),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_02152_)
  );
  OAI21X1 _08381_ (
    .A(_02795_),
    .B(_02152_),
    .C(_02151_),
    .Y(_01761_)
  );
  NOR2X1 _08382_ (
    .A(_02678_),
    .B(_02795_),
    .Y(_02153_)
  );
  AOI22X1 _08383_ (
    .A( execution_unit_0.alu_0.status_3_ ),
    .B(_02146_),
    .C(_02153_),
    .D(_02540_),
    .Y(_02154_)
  );
  NAND3X1 _08384_ (
    .A(_02540_),
    .B( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .C( execution_unit_0.alu_0.alu_stat_3_ ),
    .Y(_02155_)
  );
  OAI21X1 _08385_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .B(_02154_),
    .C(_02155_),
    .Y(_01762_)
  );
  AND2X1 _08386_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_15_ ),
    .Y(_02156_)
  );
  INVX1 _08387_ (
    .A(_02156_),
    .Y(_02157_)
  );
  NAND2X1 _08388_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02569_),
    .Y(_02158_)
  );
  NOR2X1 _08389_ (
    .A(_02156_),
    .B(_02158_),
    .Y(_02159_)
  );
  OR2X1 _08390_ (
    .A(_02156_),
    .B(_02158_),
    .Y(_02160_)
  );
  OAI21X1 _08391_ (
    .A( execution_unit_0.reg_sr_clr ),
    .B(_02541_),
    .C( execution_unit_0.alu_0.inst_bw ),
    .Y(_02161_)
  );
  INVX1 _08392_ (
    .A(_02161_),
    .Y(_02162_)
  );
  NAND2X1 _08393_ (
    .A(_02814_),
    .B(_02162_),
    .Y(_02163_)
  );
  OAI21X1 _08394_ (
    .A(_02544_),
    .B(_02566_),
    .C( execution_unit_0.reg_src_0_ ),
    .Y(_02164_)
  );
  NAND2X1 _08395_ (
    .A(_02163_),
    .B(_02164_),
    .Y(_02165_)
  );
  AOI21X1 _08396_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02569_),
    .C(_02156_),
    .Y(_02166_)
  );
  AOI22X1 _08397_ (
    .A(_02159_),
    .B(_02165_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_0_ ),
    .Y(_02167_)
  );
  OAI21X1 _08398_ (
    .A(_02551_),
    .B(_02157_),
    .C(_02167_),
    .Y(_01763_)
  );
  AOI22X1 _08399_ (
    .A(_02828_),
    .B(_02841_),
    .C(_02162_),
    .D(_02814_),
    .Y(_02168_)
  );
  OAI21X1 _08400_ (
    .A( execution_unit_0.reg_src_0_ ),
    .B(_02161_),
    .C( execution_unit_0.reg_src_1_ ),
    .Y(_02169_)
  );
  XNOR2X1 _08401_ (
    .A( execution_unit_0.reg_src_1_ ),
    .B(_02163_),
    .Y(_02170_)
  );
  AOI22X1 _08402_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_1_ ),
    .Y(_02171_)
  );
  OAI21X1 _08403_ (
    .A(_02160_),
    .B(_02170_),
    .C(_02171_),
    .Y(_01764_)
  );
  XNOR2X1 _08404_ (
    .A( execution_unit_0.reg_src_2_ ),
    .B(_02168_),
    .Y(_02172_)
  );
  AOI22X1 _08405_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_2_ ),
    .Y(_02173_)
  );
  OAI21X1 _08406_ (
    .A(_02160_),
    .B(_02172_),
    .C(_02173_),
    .Y(_01765_)
  );
  NOR3X1 _08407_ (
    .A(_02597_),
    .B(_02613_),
    .C(_02169_),
    .Y(_02174_)
  );
  NAND3X1 _08408_ (
    .A( execution_unit_0.reg_src_3_ ),
    .B( execution_unit_0.reg_src_2_ ),
    .C(_02168_),
    .Y(_02175_)
  );
  OAI21X1 _08409_ (
    .A(_02613_),
    .B(_02169_),
    .C(_02597_),
    .Y(_02176_)
  );
  NAND2X1 _08410_ (
    .A(_02175_),
    .B(_02176_),
    .Y(_02177_)
  );
  AOI22X1 _08411_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_3_ ),
    .Y(_02178_)
  );
  OAI21X1 _08412_ (
    .A(_02160_),
    .B(_02177_),
    .C(_02178_),
    .Y(_01766_)
  );
  XNOR2X1 _08413_ (
    .A(_02629_),
    .B(_02174_),
    .Y(_02179_)
  );
  AOI22X1 _08414_ (
    .A( execution_unit_0.register_file_0.r15_4_ ),
    .B(_02166_),
    .C(_02179_),
    .D(_02159_),
    .Y(_02180_)
  );
  OAI21X1 _08415_ (
    .A(_02559_),
    .B(_02157_),
    .C(_02180_),
    .Y(_01767_)
  );
  NOR3X1 _08416_ (
    .A(_02629_),
    .B(_02647_),
    .C(_02175_),
    .Y(_02181_)
  );
  NAND3X1 _08417_ (
    .A( execution_unit_0.reg_src_4_ ),
    .B( execution_unit_0.reg_src_5_ ),
    .C(_02174_),
    .Y(_02182_)
  );
  OAI21X1 _08418_ (
    .A(_02629_),
    .B(_02175_),
    .C(_02647_),
    .Y(_02183_)
  );
  NAND2X1 _08419_ (
    .A(_02182_),
    .B(_02183_),
    .Y(_02184_)
  );
  AOI22X1 _08420_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_5_ ),
    .Y(_02185_)
  );
  OAI21X1 _08421_ (
    .A(_02160_),
    .B(_02184_),
    .C(_02185_),
    .Y(_01768_)
  );
  XNOR2X1 _08422_ (
    .A(_02662_),
    .B(_02181_),
    .Y(_02186_)
  );
  AOI22X1 _08423_ (
    .A( execution_unit_0.register_file_0.r15_6_ ),
    .B(_02166_),
    .C(_02186_),
    .D(_02159_),
    .Y(_02187_)
  );
  OAI21X1 _08424_ (
    .A(_02562_),
    .B(_02157_),
    .C(_02187_),
    .Y(_01769_)
  );
  NOR3X1 _08425_ (
    .A(_02662_),
    .B(_02677_),
    .C(_02182_),
    .Y(_02188_)
  );
  NAND3X1 _08426_ (
    .A( execution_unit_0.reg_src_6_ ),
    .B( execution_unit_0.reg_src_7_ ),
    .C(_02181_),
    .Y(_02189_)
  );
  OAI21X1 _08427_ (
    .A(_02662_),
    .B(_02182_),
    .C(_02677_),
    .Y(_02190_)
  );
  NAND2X1 _08428_ (
    .A(_02189_),
    .B(_02190_),
    .Y(_02191_)
  );
  AOI22X1 _08429_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_7_ ),
    .Y(_02192_)
  );
  OAI21X1 _08430_ (
    .A(_02160_),
    .B(_02191_),
    .C(_02192_),
    .Y(_01770_)
  );
  XNOR2X1 _08431_ (
    .A( execution_unit_0.reg_src_8_ ),
    .B(_02188_),
    .Y(_02193_)
  );
  AOI22X1 _08432_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_8_ ),
    .Y(_02194_)
  );
  OAI21X1 _08433_ (
    .A(_02160_),
    .B(_02193_),
    .C(_02194_),
    .Y(_01771_)
  );
  NOR3X1 _08434_ (
    .A(_02693_),
    .B(_02708_),
    .C(_02189_),
    .Y(_02195_)
  );
  NAND3X1 _08435_ (
    .A( execution_unit_0.reg_src_8_ ),
    .B( execution_unit_0.reg_src_9_ ),
    .C(_02188_),
    .Y(_02196_)
  );
  OAI21X1 _08436_ (
    .A(_02693_),
    .B(_02189_),
    .C(_02708_),
    .Y(_02197_)
  );
  NAND2X1 _08437_ (
    .A(_02196_),
    .B(_02197_),
    .Y(_02198_)
  );
  AOI22X1 _08438_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_9_ ),
    .Y(_02199_)
  );
  OAI21X1 _08439_ (
    .A(_02160_),
    .B(_02198_),
    .C(_02199_),
    .Y(_01772_)
  );
  XNOR2X1 _08440_ (
    .A( execution_unit_0.reg_src_10_ ),
    .B(_02195_),
    .Y(_02200_)
  );
  AOI22X1 _08441_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_10_ ),
    .Y(_02201_)
  );
  OAI21X1 _08442_ (
    .A(_02160_),
    .B(_02200_),
    .C(_02201_),
    .Y(_01773_)
  );
  NOR3X1 _08443_ (
    .A(_02724_),
    .B(_02738_),
    .C(_02196_),
    .Y(_02202_)
  );
  NAND3X1 _08444_ (
    .A( execution_unit_0.reg_src_10_ ),
    .B( execution_unit_0.reg_src_11_ ),
    .C(_02195_),
    .Y(_02203_)
  );
  OAI21X1 _08445_ (
    .A(_02724_),
    .B(_02196_),
    .C(_02738_),
    .Y(_02204_)
  );
  NAND2X1 _08446_ (
    .A(_02203_),
    .B(_02204_),
    .Y(_02205_)
  );
  AOI22X1 _08447_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_11_ ),
    .Y(_02206_)
  );
  OAI21X1 _08448_ (
    .A(_02160_),
    .B(_02205_),
    .C(_02206_),
    .Y(_01774_)
  );
  XNOR2X1 _08449_ (
    .A(_02752_),
    .B(_02202_),
    .Y(_02207_)
  );
  AOI22X1 _08450_ (
    .A( execution_unit_0.register_file_0.r15_12_ ),
    .B(_02166_),
    .C(_02207_),
    .D(_02159_),
    .Y(_02208_)
  );
  OAI21X1 _08451_ (
    .A(_02739_),
    .B(_02157_),
    .C(_02208_),
    .Y(_01775_)
  );
  NOR3X1 _08452_ (
    .A(_02752_),
    .B(_02766_),
    .C(_02203_),
    .Y(_02209_)
  );
  NAND3X1 _08453_ (
    .A( execution_unit_0.reg_src_12_ ),
    .B( execution_unit_0.reg_src_13_ ),
    .C(_02202_),
    .Y(_02210_)
  );
  OAI21X1 _08454_ (
    .A(_02752_),
    .B(_02203_),
    .C(_02766_),
    .Y(_02211_)
  );
  NAND2X1 _08455_ (
    .A(_02210_),
    .B(_02211_),
    .Y(_02212_)
  );
  AOI22X1 _08456_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_13_ ),
    .Y(_02213_)
  );
  OAI21X1 _08457_ (
    .A(_02160_),
    .B(_02212_),
    .C(_02213_),
    .Y(_01776_)
  );
  XNOR2X1 _08458_ (
    .A(_02781_),
    .B(_02209_),
    .Y(_02214_)
  );
  AOI22X1 _08459_ (
    .A( execution_unit_0.register_file_0.r15_14_ ),
    .B(_02166_),
    .C(_02214_),
    .D(_02159_),
    .Y(_02215_)
  );
  OAI21X1 _08460_ (
    .A(_02767_),
    .B(_02157_),
    .C(_02215_),
    .Y(_01777_)
  );
  OAI21X1 _08461_ (
    .A(_02781_),
    .B(_02210_),
    .C(_02794_),
    .Y(_02216_)
  );
  NAND3X1 _08462_ (
    .A( execution_unit_0.reg_src_14_ ),
    .B( execution_unit_0.reg_src_15_ ),
    .C(_02209_),
    .Y(_02217_)
  );
  NAND2X1 _08463_ (
    .A(_02216_),
    .B(_02217_),
    .Y(_02218_)
  );
  AOI22X1 _08464_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02156_),
    .C(_02166_),
    .D( execution_unit_0.register_file_0.r15_15_ ),
    .Y(_02219_)
  );
  OAI21X1 _08465_ (
    .A(_02160_),
    .B(_02218_),
    .C(_02219_),
    .Y(_01778_)
  );
  AND2X1 _08466_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_14_ ),
    .Y(_02220_)
  );
  NAND2X1 _08467_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_14_ ),
    .Y(_02221_)
  );
  NAND2X1 _08468_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02580_),
    .Y(_02222_)
  );
  NOR2X1 _08469_ (
    .A(_02220_),
    .B(_02222_),
    .Y(_02223_)
  );
  OR2X1 _08470_ (
    .A(_02220_),
    .B(_02222_),
    .Y(_02224_)
  );
  AOI21X1 _08471_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02580_),
    .C(_02220_),
    .Y(_02225_)
  );
  INVX1 _08472_ (
    .A(_02225_),
    .Y(_02226_)
  );
  OAI22X1 _08473_ (
    .A(_02165_),
    .B(_02224_),
    .C(_02226_),
    .D( execution_unit_0.register_file_0.r14_0_ ),
    .Y(_02227_)
  );
  AOI21X1 _08474_ (
    .A(_02551_),
    .B(_02220_),
    .C(_02227_),
    .Y(_01779_)
  );
  AOI22X1 _08475_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_1_ ),
    .Y(_02228_)
  );
  OAI21X1 _08476_ (
    .A(_02170_),
    .B(_02224_),
    .C(_02228_),
    .Y(_01780_)
  );
  AOI22X1 _08477_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_2_ ),
    .Y(_02229_)
  );
  OAI21X1 _08478_ (
    .A(_02172_),
    .B(_02224_),
    .C(_02229_),
    .Y(_01781_)
  );
  AOI22X1 _08479_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_3_ ),
    .Y(_02230_)
  );
  OAI21X1 _08480_ (
    .A(_02177_),
    .B(_02224_),
    .C(_02230_),
    .Y(_01782_)
  );
  AOI22X1 _08481_ (
    .A(_02179_),
    .B(_02223_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_4_ ),
    .Y(_02231_)
  );
  OAI21X1 _08482_ (
    .A(_02559_),
    .B(_02221_),
    .C(_02231_),
    .Y(_01783_)
  );
  AOI22X1 _08483_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_5_ ),
    .Y(_02232_)
  );
  OAI21X1 _08484_ (
    .A(_02184_),
    .B(_02224_),
    .C(_02232_),
    .Y(_01784_)
  );
  AOI22X1 _08485_ (
    .A(_02186_),
    .B(_02223_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_6_ ),
    .Y(_02233_)
  );
  OAI21X1 _08486_ (
    .A(_02562_),
    .B(_02221_),
    .C(_02233_),
    .Y(_01785_)
  );
  AOI22X1 _08487_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_7_ ),
    .Y(_02234_)
  );
  OAI21X1 _08488_ (
    .A(_02191_),
    .B(_02224_),
    .C(_02234_),
    .Y(_01786_)
  );
  AOI22X1 _08489_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_8_ ),
    .Y(_02235_)
  );
  OAI21X1 _08490_ (
    .A(_02193_),
    .B(_02224_),
    .C(_02235_),
    .Y(_01787_)
  );
  AOI22X1 _08491_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_9_ ),
    .Y(_02236_)
  );
  OAI21X1 _08492_ (
    .A(_02198_),
    .B(_02224_),
    .C(_02236_),
    .Y(_01788_)
  );
  AOI22X1 _08493_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_10_ ),
    .Y(_02237_)
  );
  OAI21X1 _08494_ (
    .A(_02200_),
    .B(_02224_),
    .C(_02237_),
    .Y(_01789_)
  );
  AOI22X1 _08495_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_11_ ),
    .Y(_02238_)
  );
  OAI21X1 _08496_ (
    .A(_02205_),
    .B(_02224_),
    .C(_02238_),
    .Y(_01790_)
  );
  AOI22X1 _08497_ (
    .A(_02207_),
    .B(_02223_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_12_ ),
    .Y(_02239_)
  );
  OAI21X1 _08498_ (
    .A(_02739_),
    .B(_02221_),
    .C(_02239_),
    .Y(_01791_)
  );
  AOI22X1 _08499_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_13_ ),
    .Y(_02240_)
  );
  OAI21X1 _08500_ (
    .A(_02212_),
    .B(_02224_),
    .C(_02240_),
    .Y(_01792_)
  );
  AOI22X1 _08501_ (
    .A(_02214_),
    .B(_02223_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_14_ ),
    .Y(_02241_)
  );
  OAI21X1 _08502_ (
    .A(_02767_),
    .B(_02221_),
    .C(_02241_),
    .Y(_01793_)
  );
  AOI22X1 _08503_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02220_),
    .C(_02225_),
    .D( execution_unit_0.register_file_0.r14_15_ ),
    .Y(_02242_)
  );
  OAI21X1 _08504_ (
    .A(_02218_),
    .B(_02224_),
    .C(_02242_),
    .Y(_01794_)
  );
  AND2X1 _08505_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_13_ ),
    .Y(_02243_)
  );
  NAND2X1 _08506_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_13_ ),
    .Y(_02244_)
  );
  NAND2X1 _08507_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02568_),
    .Y(_02245_)
  );
  NOR2X1 _08508_ (
    .A(_02243_),
    .B(_02245_),
    .Y(_02246_)
  );
  OR2X1 _08509_ (
    .A(_02243_),
    .B(_02245_),
    .Y(_02247_)
  );
  AOI21X1 _08510_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02568_),
    .C(_02243_),
    .Y(_02248_)
  );
  INVX1 _08511_ (
    .A(_02248_),
    .Y(_02249_)
  );
  OAI22X1 _08512_ (
    .A(_02165_),
    .B(_02247_),
    .C(_02249_),
    .D( execution_unit_0.register_file_0.r13_0_ ),
    .Y(_02250_)
  );
  AOI21X1 _08513_ (
    .A(_02551_),
    .B(_02243_),
    .C(_02250_),
    .Y(_01795_)
  );
  AOI22X1 _08514_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_1_ ),
    .Y(_02251_)
  );
  OAI21X1 _08515_ (
    .A(_02170_),
    .B(_02247_),
    .C(_02251_),
    .Y(_01796_)
  );
  AOI22X1 _08516_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_2_ ),
    .Y(_02252_)
  );
  OAI21X1 _08517_ (
    .A(_02172_),
    .B(_02247_),
    .C(_02252_),
    .Y(_01797_)
  );
  AOI22X1 _08518_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_3_ ),
    .Y(_02253_)
  );
  OAI21X1 _08519_ (
    .A(_02177_),
    .B(_02247_),
    .C(_02253_),
    .Y(_01798_)
  );
  AOI22X1 _08520_ (
    .A(_02179_),
    .B(_02246_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_4_ ),
    .Y(_02254_)
  );
  OAI21X1 _08521_ (
    .A(_02559_),
    .B(_02244_),
    .C(_02254_),
    .Y(_01799_)
  );
  AOI22X1 _08522_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_5_ ),
    .Y(_02255_)
  );
  OAI21X1 _08523_ (
    .A(_02184_),
    .B(_02247_),
    .C(_02255_),
    .Y(_01800_)
  );
  AOI22X1 _08524_ (
    .A(_02186_),
    .B(_02246_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_6_ ),
    .Y(_02256_)
  );
  OAI21X1 _08525_ (
    .A(_02562_),
    .B(_02244_),
    .C(_02256_),
    .Y(_01801_)
  );
  AOI22X1 _08526_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_7_ ),
    .Y(_02257_)
  );
  OAI21X1 _08527_ (
    .A(_02191_),
    .B(_02247_),
    .C(_02257_),
    .Y(_01802_)
  );
  AOI22X1 _08528_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_8_ ),
    .Y(_02258_)
  );
  OAI21X1 _08529_ (
    .A(_02193_),
    .B(_02247_),
    .C(_02258_),
    .Y(_01803_)
  );
  AOI22X1 _08530_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_9_ ),
    .Y(_02259_)
  );
  OAI21X1 _08531_ (
    .A(_02198_),
    .B(_02247_),
    .C(_02259_),
    .Y(_01804_)
  );
  AOI22X1 _08532_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_10_ ),
    .Y(_02260_)
  );
  OAI21X1 _08533_ (
    .A(_02200_),
    .B(_02247_),
    .C(_02260_),
    .Y(_01805_)
  );
  AOI22X1 _08534_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_11_ ),
    .Y(_02261_)
  );
  OAI21X1 _08535_ (
    .A(_02205_),
    .B(_02247_),
    .C(_02261_),
    .Y(_01806_)
  );
  AOI22X1 _08536_ (
    .A(_02207_),
    .B(_02246_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_12_ ),
    .Y(_02262_)
  );
  OAI21X1 _08537_ (
    .A(_02739_),
    .B(_02244_),
    .C(_02262_),
    .Y(_01807_)
  );
  AOI22X1 _08538_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_13_ ),
    .Y(_02263_)
  );
  OAI21X1 _08539_ (
    .A(_02212_),
    .B(_02247_),
    .C(_02263_),
    .Y(_01808_)
  );
  AOI22X1 _08540_ (
    .A(_02214_),
    .B(_02246_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_14_ ),
    .Y(_02264_)
  );
  OAI21X1 _08541_ (
    .A(_02767_),
    .B(_02244_),
    .C(_02264_),
    .Y(_01809_)
  );
  AOI22X1 _08542_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02243_),
    .C(_02248_),
    .D( execution_unit_0.register_file_0.r13_15_ ),
    .Y(_02265_)
  );
  OAI21X1 _08543_ (
    .A(_02218_),
    .B(_02247_),
    .C(_02265_),
    .Y(_01810_)
  );
  AND2X1 _08544_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_12_ ),
    .Y(_02266_)
  );
  NAND2X1 _08545_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_12_ ),
    .Y(_02267_)
  );
  NAND2X1 _08546_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02593_),
    .Y(_02268_)
  );
  NOR2X1 _08547_ (
    .A(_02266_),
    .B(_02268_),
    .Y(_02269_)
  );
  OR2X1 _08548_ (
    .A(_02266_),
    .B(_02268_),
    .Y(_02270_)
  );
  AOI21X1 _08549_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02593_),
    .C(_02266_),
    .Y(_02271_)
  );
  INVX1 _08550_ (
    .A(_02271_),
    .Y(_02272_)
  );
  OAI22X1 _08551_ (
    .A(_02165_),
    .B(_02270_),
    .C(_02272_),
    .D( execution_unit_0.register_file_0.r12_0_ ),
    .Y(_02273_)
  );
  AOI21X1 _08552_ (
    .A(_02551_),
    .B(_02266_),
    .C(_02273_),
    .Y(_01811_)
  );
  AOI22X1 _08553_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_1_ ),
    .Y(_02274_)
  );
  OAI21X1 _08554_ (
    .A(_02170_),
    .B(_02270_),
    .C(_02274_),
    .Y(_01812_)
  );
  AOI22X1 _08555_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_2_ ),
    .Y(_02275_)
  );
  OAI21X1 _08556_ (
    .A(_02172_),
    .B(_02270_),
    .C(_02275_),
    .Y(_01813_)
  );
  AOI22X1 _08557_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_3_ ),
    .Y(_02276_)
  );
  OAI21X1 _08558_ (
    .A(_02177_),
    .B(_02270_),
    .C(_02276_),
    .Y(_01814_)
  );
  AOI22X1 _08559_ (
    .A(_02179_),
    .B(_02269_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_4_ ),
    .Y(_02277_)
  );
  OAI21X1 _08560_ (
    .A(_02559_),
    .B(_02267_),
    .C(_02277_),
    .Y(_01815_)
  );
  AOI22X1 _08561_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_5_ ),
    .Y(_02278_)
  );
  OAI21X1 _08562_ (
    .A(_02184_),
    .B(_02270_),
    .C(_02278_),
    .Y(_01816_)
  );
  AOI22X1 _08563_ (
    .A(_02186_),
    .B(_02269_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_6_ ),
    .Y(_02279_)
  );
  OAI21X1 _08564_ (
    .A(_02562_),
    .B(_02267_),
    .C(_02279_),
    .Y(_01817_)
  );
  AOI22X1 _08565_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_7_ ),
    .Y(_02280_)
  );
  OAI21X1 _08566_ (
    .A(_02191_),
    .B(_02270_),
    .C(_02280_),
    .Y(_01818_)
  );
  AOI22X1 _08567_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_8_ ),
    .Y(_02281_)
  );
  OAI21X1 _08568_ (
    .A(_02193_),
    .B(_02270_),
    .C(_02281_),
    .Y(_01819_)
  );
  AOI22X1 _08569_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_9_ ),
    .Y(_02282_)
  );
  OAI21X1 _08570_ (
    .A(_02198_),
    .B(_02270_),
    .C(_02282_),
    .Y(_01820_)
  );
  AOI22X1 _08571_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_10_ ),
    .Y(_02283_)
  );
  OAI21X1 _08572_ (
    .A(_02200_),
    .B(_02270_),
    .C(_02283_),
    .Y(_01821_)
  );
  AOI22X1 _08573_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_11_ ),
    .Y(_02284_)
  );
  OAI21X1 _08574_ (
    .A(_02205_),
    .B(_02270_),
    .C(_02284_),
    .Y(_01822_)
  );
  AOI22X1 _08575_ (
    .A(_02207_),
    .B(_02269_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_12_ ),
    .Y(_02285_)
  );
  OAI21X1 _08576_ (
    .A(_02739_),
    .B(_02267_),
    .C(_02285_),
    .Y(_01823_)
  );
  AOI22X1 _08577_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_13_ ),
    .Y(_02286_)
  );
  OAI21X1 _08578_ (
    .A(_02212_),
    .B(_02270_),
    .C(_02286_),
    .Y(_01824_)
  );
  AOI22X1 _08579_ (
    .A(_02214_),
    .B(_02269_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_14_ ),
    .Y(_02287_)
  );
  OAI21X1 _08580_ (
    .A(_02767_),
    .B(_02267_),
    .C(_02287_),
    .Y(_01825_)
  );
  AOI22X1 _08581_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02266_),
    .C(_02271_),
    .D( execution_unit_0.register_file_0.r12_15_ ),
    .Y(_02288_)
  );
  OAI21X1 _08582_ (
    .A(_02218_),
    .B(_02270_),
    .C(_02288_),
    .Y(_01826_)
  );
  AND2X1 _08583_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_11_ ),
    .Y(_02289_)
  );
  NAND2X1 _08584_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_11_ ),
    .Y(_02290_)
  );
  NAND2X1 _08585_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02591_),
    .Y(_02291_)
  );
  NOR2X1 _08586_ (
    .A(_02289_),
    .B(_02291_),
    .Y(_02292_)
  );
  OR2X1 _08587_ (
    .A(_02289_),
    .B(_02291_),
    .Y(_02293_)
  );
  AOI21X1 _08588_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02591_),
    .C(_02289_),
    .Y(_02294_)
  );
  NAND2X1 _08589_ (
    .A(_02550_),
    .B(_02294_),
    .Y(_02295_)
  );
  OAI21X1 _08590_ (
    .A(_02165_),
    .B(_02293_),
    .C(_02295_),
    .Y(_02296_)
  );
  AOI21X1 _08591_ (
    .A(_02551_),
    .B(_02289_),
    .C(_02296_),
    .Y(_01827_)
  );
  AOI22X1 _08592_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_1_ ),
    .Y(_02297_)
  );
  OAI21X1 _08593_ (
    .A(_02170_),
    .B(_02293_),
    .C(_02297_),
    .Y(_01828_)
  );
  AOI22X1 _08594_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_2_ ),
    .Y(_02298_)
  );
  OAI21X1 _08595_ (
    .A(_02172_),
    .B(_02293_),
    .C(_02298_),
    .Y(_01829_)
  );
  AOI22X1 _08596_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_3_ ),
    .Y(_02299_)
  );
  OAI21X1 _08597_ (
    .A(_02177_),
    .B(_02293_),
    .C(_02299_),
    .Y(_01830_)
  );
  AOI22X1 _08598_ (
    .A(_02179_),
    .B(_02292_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_4_ ),
    .Y(_02300_)
  );
  OAI21X1 _08599_ (
    .A(_02559_),
    .B(_02290_),
    .C(_02300_),
    .Y(_01831_)
  );
  AOI22X1 _08600_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_5_ ),
    .Y(_02301_)
  );
  OAI21X1 _08601_ (
    .A(_02184_),
    .B(_02293_),
    .C(_02301_),
    .Y(_01832_)
  );
  AOI22X1 _08602_ (
    .A(_02186_),
    .B(_02292_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_6_ ),
    .Y(_02302_)
  );
  OAI21X1 _08603_ (
    .A(_02562_),
    .B(_02290_),
    .C(_02302_),
    .Y(_01833_)
  );
  AOI22X1 _08604_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_7_ ),
    .Y(_02303_)
  );
  OAI21X1 _08605_ (
    .A(_02191_),
    .B(_02293_),
    .C(_02303_),
    .Y(_01834_)
  );
  AOI22X1 _08606_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_8_ ),
    .Y(_02304_)
  );
  OAI21X1 _08607_ (
    .A(_02193_),
    .B(_02293_),
    .C(_02304_),
    .Y(_01835_)
  );
  AOI22X1 _08608_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_9_ ),
    .Y(_02305_)
  );
  OAI21X1 _08609_ (
    .A(_02198_),
    .B(_02293_),
    .C(_02305_),
    .Y(_01836_)
  );
  AOI22X1 _08610_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_10_ ),
    .Y(_02306_)
  );
  OAI21X1 _08611_ (
    .A(_02200_),
    .B(_02293_),
    .C(_02306_),
    .Y(_01837_)
  );
  AOI22X1 _08612_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_11_ ),
    .Y(_02307_)
  );
  OAI21X1 _08613_ (
    .A(_02205_),
    .B(_02293_),
    .C(_02307_),
    .Y(_01838_)
  );
  AOI22X1 _08614_ (
    .A(_02207_),
    .B(_02292_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_12_ ),
    .Y(_02308_)
  );
  OAI21X1 _08615_ (
    .A(_02739_),
    .B(_02290_),
    .C(_02308_),
    .Y(_01839_)
  );
  AOI22X1 _08616_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_13_ ),
    .Y(_02309_)
  );
  OAI21X1 _08617_ (
    .A(_02212_),
    .B(_02293_),
    .C(_02309_),
    .Y(_01840_)
  );
  AOI22X1 _08618_ (
    .A(_02214_),
    .B(_02292_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_14_ ),
    .Y(_02310_)
  );
  OAI21X1 _08619_ (
    .A(_02767_),
    .B(_02290_),
    .C(_02310_),
    .Y(_01841_)
  );
  AOI22X1 _08620_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02289_),
    .C(_02294_),
    .D( execution_unit_0.register_file_0.r11_15_ ),
    .Y(_02311_)
  );
  OAI21X1 _08621_ (
    .A(_02218_),
    .B(_02293_),
    .C(_02311_),
    .Y(_01842_)
  );
  AND2X1 _08622_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_10_ ),
    .Y(_02312_)
  );
  NAND2X1 _08623_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_10_ ),
    .Y(_02313_)
  );
  NAND2X1 _08624_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02583_),
    .Y(_02314_)
  );
  NOR2X1 _08625_ (
    .A(_02312_),
    .B(_02314_),
    .Y(_02315_)
  );
  OR2X1 _08626_ (
    .A(_02312_),
    .B(_02314_),
    .Y(_02316_)
  );
  AOI21X1 _08627_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02583_),
    .C(_02312_),
    .Y(_02317_)
  );
  NAND2X1 _08628_ (
    .A(_02549_),
    .B(_02317_),
    .Y(_02318_)
  );
  OAI21X1 _08629_ (
    .A(_02165_),
    .B(_02316_),
    .C(_02318_),
    .Y(_02319_)
  );
  AOI21X1 _08630_ (
    .A(_02551_),
    .B(_02312_),
    .C(_02319_),
    .Y(_01843_)
  );
  AOI22X1 _08631_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_1_ ),
    .Y(_02320_)
  );
  OAI21X1 _08632_ (
    .A(_02170_),
    .B(_02316_),
    .C(_02320_),
    .Y(_01844_)
  );
  AOI22X1 _08633_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_2_ ),
    .Y(_02321_)
  );
  OAI21X1 _08634_ (
    .A(_02172_),
    .B(_02316_),
    .C(_02321_),
    .Y(_01845_)
  );
  AOI22X1 _08635_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_3_ ),
    .Y(_02322_)
  );
  OAI21X1 _08636_ (
    .A(_02177_),
    .B(_02316_),
    .C(_02322_),
    .Y(_01846_)
  );
  AOI22X1 _08637_ (
    .A(_02179_),
    .B(_02315_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_4_ ),
    .Y(_02323_)
  );
  OAI21X1 _08638_ (
    .A(_02559_),
    .B(_02313_),
    .C(_02323_),
    .Y(_01847_)
  );
  AOI22X1 _08639_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_5_ ),
    .Y(_02324_)
  );
  OAI21X1 _08640_ (
    .A(_02184_),
    .B(_02316_),
    .C(_02324_),
    .Y(_01848_)
  );
  AOI22X1 _08641_ (
    .A(_02186_),
    .B(_02315_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_6_ ),
    .Y(_02325_)
  );
  OAI21X1 _08642_ (
    .A(_02562_),
    .B(_02313_),
    .C(_02325_),
    .Y(_01849_)
  );
  AOI22X1 _08643_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_7_ ),
    .Y(_02326_)
  );
  OAI21X1 _08644_ (
    .A(_02191_),
    .B(_02316_),
    .C(_02326_),
    .Y(_01850_)
  );
  AOI22X1 _08645_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_8_ ),
    .Y(_02327_)
  );
  OAI21X1 _08646_ (
    .A(_02193_),
    .B(_02316_),
    .C(_02327_),
    .Y(_01851_)
  );
  AOI22X1 _08647_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_9_ ),
    .Y(_02328_)
  );
  OAI21X1 _08648_ (
    .A(_02198_),
    .B(_02316_),
    .C(_02328_),
    .Y(_01852_)
  );
  AOI22X1 _08649_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_10_ ),
    .Y(_02329_)
  );
  OAI21X1 _08650_ (
    .A(_02200_),
    .B(_02316_),
    .C(_02329_),
    .Y(_01853_)
  );
  AOI22X1 _08651_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_11_ ),
    .Y(_02330_)
  );
  OAI21X1 _08652_ (
    .A(_02205_),
    .B(_02316_),
    .C(_02330_),
    .Y(_01854_)
  );
  AOI22X1 _08653_ (
    .A(_02207_),
    .B(_02315_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_12_ ),
    .Y(_02331_)
  );
  OAI21X1 _08654_ (
    .A(_02739_),
    .B(_02313_),
    .C(_02331_),
    .Y(_01855_)
  );
  AOI22X1 _08655_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_13_ ),
    .Y(_02332_)
  );
  OAI21X1 _08656_ (
    .A(_02212_),
    .B(_02316_),
    .C(_02332_),
    .Y(_01856_)
  );
  AOI22X1 _08657_ (
    .A(_02214_),
    .B(_02315_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_14_ ),
    .Y(_02333_)
  );
  OAI21X1 _08658_ (
    .A(_02767_),
    .B(_02313_),
    .C(_02333_),
    .Y(_01857_)
  );
  AOI22X1 _08659_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02312_),
    .C(_02317_),
    .D( execution_unit_0.register_file_0.r10_15_ ),
    .Y(_02334_)
  );
  OAI21X1 _08660_ (
    .A(_02218_),
    .B(_02316_),
    .C(_02334_),
    .Y(_01858_)
  );
  AND2X1 _08661_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_9_ ),
    .Y(_02335_)
  );
  NAND2X1 _08662_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_9_ ),
    .Y(_02336_)
  );
  NAND2X1 _08663_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02588_),
    .Y(_02337_)
  );
  NOR2X1 _08664_ (
    .A(_02335_),
    .B(_02337_),
    .Y(_02338_)
  );
  OR2X1 _08665_ (
    .A(_02335_),
    .B(_02337_),
    .Y(_02339_)
  );
  AOI21X1 _08666_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02588_),
    .C(_02335_),
    .Y(_02340_)
  );
  INVX1 _08667_ (
    .A(_02340_),
    .Y(_02341_)
  );
  OAI22X1 _08668_ (
    .A(_02165_),
    .B(_02339_),
    .C(_02341_),
    .D( execution_unit_0.register_file_0.r9_0_ ),
    .Y(_02342_)
  );
  AOI21X1 _08669_ (
    .A(_02551_),
    .B(_02335_),
    .C(_02342_),
    .Y(_01859_)
  );
  AOI22X1 _08670_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_1_ ),
    .Y(_02343_)
  );
  OAI21X1 _08671_ (
    .A(_02170_),
    .B(_02339_),
    .C(_02343_),
    .Y(_01860_)
  );
  AOI22X1 _08672_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_2_ ),
    .Y(_02344_)
  );
  OAI21X1 _08673_ (
    .A(_02172_),
    .B(_02339_),
    .C(_02344_),
    .Y(_01861_)
  );
  AOI22X1 _08674_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_3_ ),
    .Y(_02345_)
  );
  OAI21X1 _08675_ (
    .A(_02177_),
    .B(_02339_),
    .C(_02345_),
    .Y(_01862_)
  );
  AOI22X1 _08676_ (
    .A(_02179_),
    .B(_02338_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_4_ ),
    .Y(_02346_)
  );
  OAI21X1 _08677_ (
    .A(_02559_),
    .B(_02336_),
    .C(_02346_),
    .Y(_01863_)
  );
  AOI22X1 _08678_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_5_ ),
    .Y(_02347_)
  );
  OAI21X1 _08679_ (
    .A(_02184_),
    .B(_02339_),
    .C(_02347_),
    .Y(_01864_)
  );
  AOI22X1 _08680_ (
    .A(_02186_),
    .B(_02338_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_6_ ),
    .Y(_02348_)
  );
  OAI21X1 _08681_ (
    .A(_02562_),
    .B(_02336_),
    .C(_02348_),
    .Y(_01865_)
  );
  AOI22X1 _08682_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_7_ ),
    .Y(_02349_)
  );
  OAI21X1 _08683_ (
    .A(_02191_),
    .B(_02339_),
    .C(_02349_),
    .Y(_01866_)
  );
  AOI22X1 _08684_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_8_ ),
    .Y(_02350_)
  );
  OAI21X1 _08685_ (
    .A(_02193_),
    .B(_02339_),
    .C(_02350_),
    .Y(_01867_)
  );
  AOI22X1 _08686_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_9_ ),
    .Y(_02351_)
  );
  OAI21X1 _08687_ (
    .A(_02198_),
    .B(_02339_),
    .C(_02351_),
    .Y(_01868_)
  );
  AOI22X1 _08688_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_10_ ),
    .Y(_02352_)
  );
  OAI21X1 _08689_ (
    .A(_02200_),
    .B(_02339_),
    .C(_02352_),
    .Y(_01869_)
  );
  AOI22X1 _08690_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_11_ ),
    .Y(_02353_)
  );
  OAI21X1 _08691_ (
    .A(_02205_),
    .B(_02339_),
    .C(_02353_),
    .Y(_01870_)
  );
  AOI22X1 _08692_ (
    .A(_02207_),
    .B(_02338_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_12_ ),
    .Y(_02354_)
  );
  OAI21X1 _08693_ (
    .A(_02739_),
    .B(_02336_),
    .C(_02354_),
    .Y(_01871_)
  );
  AOI22X1 _08694_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_13_ ),
    .Y(_02355_)
  );
  OAI21X1 _08695_ (
    .A(_02212_),
    .B(_02339_),
    .C(_02355_),
    .Y(_01872_)
  );
  AOI22X1 _08696_ (
    .A(_02214_),
    .B(_02338_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_14_ ),
    .Y(_02356_)
  );
  OAI21X1 _08697_ (
    .A(_02767_),
    .B(_02336_),
    .C(_02356_),
    .Y(_01873_)
  );
  AOI22X1 _08698_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02335_),
    .C(_02340_),
    .D( execution_unit_0.register_file_0.r9_15_ ),
    .Y(_02357_)
  );
  OAI21X1 _08699_ (
    .A(_02218_),
    .B(_02339_),
    .C(_02357_),
    .Y(_01874_)
  );
  AND2X1 _08700_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_8_ ),
    .Y(_02358_)
  );
  NAND2X1 _08701_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_8_ ),
    .Y(_02359_)
  );
  NAND2X1 _08702_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02581_),
    .Y(_02360_)
  );
  NOR2X1 _08703_ (
    .A(_02358_),
    .B(_02360_),
    .Y(_02361_)
  );
  OR2X1 _08704_ (
    .A(_02358_),
    .B(_02360_),
    .Y(_02362_)
  );
  AOI21X1 _08705_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02581_),
    .C(_02358_),
    .Y(_02363_)
  );
  OAI22X1 _08706_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02359_),
    .C(_02362_),
    .D(_02165_),
    .Y(_02364_)
  );
  AOI21X1 _08707_ (
    .A(_02548_),
    .B(_02363_),
    .C(_02364_),
    .Y(_01875_)
  );
  AOI22X1 _08708_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_1_ ),
    .Y(_02365_)
  );
  OAI21X1 _08709_ (
    .A(_02170_),
    .B(_02362_),
    .C(_02365_),
    .Y(_01876_)
  );
  AOI22X1 _08710_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_2_ ),
    .Y(_02366_)
  );
  OAI21X1 _08711_ (
    .A(_02172_),
    .B(_02362_),
    .C(_02366_),
    .Y(_01877_)
  );
  AOI22X1 _08712_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_3_ ),
    .Y(_02367_)
  );
  OAI21X1 _08713_ (
    .A(_02177_),
    .B(_02362_),
    .C(_02367_),
    .Y(_01878_)
  );
  AOI22X1 _08714_ (
    .A(_02179_),
    .B(_02361_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_4_ ),
    .Y(_02368_)
  );
  OAI21X1 _08715_ (
    .A(_02559_),
    .B(_02359_),
    .C(_02368_),
    .Y(_01879_)
  );
  AOI22X1 _08716_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_5_ ),
    .Y(_02369_)
  );
  OAI21X1 _08717_ (
    .A(_02184_),
    .B(_02362_),
    .C(_02369_),
    .Y(_01880_)
  );
  AOI22X1 _08718_ (
    .A(_02186_),
    .B(_02361_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_6_ ),
    .Y(_02370_)
  );
  OAI21X1 _08719_ (
    .A(_02562_),
    .B(_02359_),
    .C(_02370_),
    .Y(_01881_)
  );
  AOI22X1 _08720_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_7_ ),
    .Y(_02371_)
  );
  OAI21X1 _08721_ (
    .A(_02191_),
    .B(_02362_),
    .C(_02371_),
    .Y(_01882_)
  );
  AOI22X1 _08722_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_8_ ),
    .Y(_02372_)
  );
  OAI21X1 _08723_ (
    .A(_02193_),
    .B(_02362_),
    .C(_02372_),
    .Y(_01883_)
  );
  AOI22X1 _08724_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_9_ ),
    .Y(_02373_)
  );
  OAI21X1 _08725_ (
    .A(_02198_),
    .B(_02362_),
    .C(_02373_),
    .Y(_01884_)
  );
  AOI22X1 _08726_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_10_ ),
    .Y(_02374_)
  );
  OAI21X1 _08727_ (
    .A(_02200_),
    .B(_02362_),
    .C(_02374_),
    .Y(_01885_)
  );
  AOI22X1 _08728_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_11_ ),
    .Y(_02375_)
  );
  OAI21X1 _08729_ (
    .A(_02205_),
    .B(_02362_),
    .C(_02375_),
    .Y(_01886_)
  );
  AOI22X1 _08730_ (
    .A(_02207_),
    .B(_02361_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_12_ ),
    .Y(_02376_)
  );
  OAI21X1 _08731_ (
    .A(_02739_),
    .B(_02359_),
    .C(_02376_),
    .Y(_01887_)
  );
  AOI22X1 _08732_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_13_ ),
    .Y(_02377_)
  );
  OAI21X1 _08733_ (
    .A(_02212_),
    .B(_02362_),
    .C(_02377_),
    .Y(_01888_)
  );
  AOI22X1 _08734_ (
    .A(_02214_),
    .B(_02361_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_14_ ),
    .Y(_02378_)
  );
  OAI21X1 _08735_ (
    .A(_02767_),
    .B(_02359_),
    .C(_02378_),
    .Y(_01889_)
  );
  AOI22X1 _08736_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02358_),
    .C(_02363_),
    .D( execution_unit_0.register_file_0.r8_15_ ),
    .Y(_02379_)
  );
  OAI21X1 _08737_ (
    .A(_02218_),
    .B(_02362_),
    .C(_02379_),
    .Y(_01890_)
  );
  AND2X1 _08738_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_7_ ),
    .Y(_02380_)
  );
  NAND2X1 _08739_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_7_ ),
    .Y(_02381_)
  );
  NAND2X1 _08740_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02585_),
    .Y(_02382_)
  );
  NOR2X1 _08741_ (
    .A(_02380_),
    .B(_02382_),
    .Y(_02383_)
  );
  OR2X1 _08742_ (
    .A(_02380_),
    .B(_02382_),
    .Y(_02384_)
  );
  AOI21X1 _08743_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02585_),
    .C(_02380_),
    .Y(_02385_)
  );
  OAI22X1 _08744_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02381_),
    .C(_02384_),
    .D(_02165_),
    .Y(_02386_)
  );
  AOI21X1 _08745_ (
    .A(_02547_),
    .B(_02385_),
    .C(_02386_),
    .Y(_01891_)
  );
  AOI22X1 _08746_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02387_)
  );
  OAI21X1 _08747_ (
    .A(_02170_),
    .B(_02384_),
    .C(_02387_),
    .Y(_01892_)
  );
  AOI22X1 _08748_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_2_ ),
    .Y(_02388_)
  );
  OAI21X1 _08749_ (
    .A(_02172_),
    .B(_02384_),
    .C(_02388_),
    .Y(_01893_)
  );
  AOI22X1 _08750_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02389_)
  );
  OAI21X1 _08751_ (
    .A(_02177_),
    .B(_02384_),
    .C(_02389_),
    .Y(_01894_)
  );
  AOI22X1 _08752_ (
    .A(_02179_),
    .B(_02383_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_4_ ),
    .Y(_02390_)
  );
  OAI21X1 _08753_ (
    .A(_02559_),
    .B(_02381_),
    .C(_02390_),
    .Y(_01895_)
  );
  AOI22X1 _08754_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_5_ ),
    .Y(_02391_)
  );
  OAI21X1 _08755_ (
    .A(_02184_),
    .B(_02384_),
    .C(_02391_),
    .Y(_01896_)
  );
  AOI22X1 _08756_ (
    .A(_02186_),
    .B(_02383_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_6_ ),
    .Y(_02392_)
  );
  OAI21X1 _08757_ (
    .A(_02562_),
    .B(_02381_),
    .C(_02392_),
    .Y(_01897_)
  );
  AOI22X1 _08758_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_7_ ),
    .Y(_02393_)
  );
  OAI21X1 _08759_ (
    .A(_02191_),
    .B(_02384_),
    .C(_02393_),
    .Y(_01898_)
  );
  AOI22X1 _08760_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_8_ ),
    .Y(_02394_)
  );
  OAI21X1 _08761_ (
    .A(_02193_),
    .B(_02384_),
    .C(_02394_),
    .Y(_01899_)
  );
  AOI22X1 _08762_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_9_ ),
    .Y(_02395_)
  );
  OAI21X1 _08763_ (
    .A(_02198_),
    .B(_02384_),
    .C(_02395_),
    .Y(_01900_)
  );
  AOI22X1 _08764_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_10_ ),
    .Y(_02396_)
  );
  OAI21X1 _08765_ (
    .A(_02200_),
    .B(_02384_),
    .C(_02396_),
    .Y(_01901_)
  );
  AOI22X1 _08766_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_11_ ),
    .Y(_02397_)
  );
  OAI21X1 _08767_ (
    .A(_02205_),
    .B(_02384_),
    .C(_02397_),
    .Y(_01902_)
  );
  AOI22X1 _08768_ (
    .A(_02207_),
    .B(_02383_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_12_ ),
    .Y(_02398_)
  );
  OAI21X1 _08769_ (
    .A(_02739_),
    .B(_02381_),
    .C(_02398_),
    .Y(_01903_)
  );
  AOI22X1 _08770_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_13_ ),
    .Y(_02399_)
  );
  OAI21X1 _08771_ (
    .A(_02212_),
    .B(_02384_),
    .C(_02399_),
    .Y(_01904_)
  );
  AOI22X1 _08772_ (
    .A(_02214_),
    .B(_02383_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_14_ ),
    .Y(_02400_)
  );
  OAI21X1 _08773_ (
    .A(_02767_),
    .B(_02381_),
    .C(_02400_),
    .Y(_01905_)
  );
  AOI22X1 _08774_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02380_),
    .C(_02385_),
    .D( execution_unit_0.register_file_0.r7_15_ ),
    .Y(_02401_)
  );
  OAI21X1 _08775_ (
    .A(_02218_),
    .B(_02384_),
    .C(_02401_),
    .Y(_01906_)
  );
  AND2X1 _08776_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_6_ ),
    .Y(_02402_)
  );
  NAND2X1 _08777_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_6_ ),
    .Y(_02403_)
  );
  NAND2X1 _08778_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02575_),
    .Y(_02404_)
  );
  NOR2X1 _08779_ (
    .A(_02402_),
    .B(_02404_),
    .Y(_02405_)
  );
  OR2X1 _08780_ (
    .A(_02402_),
    .B(_02404_),
    .Y(_02406_)
  );
  AOI21X1 _08781_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02575_),
    .C(_02402_),
    .Y(_02407_)
  );
  OAI22X1 _08782_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02403_),
    .C(_02406_),
    .D(_02165_),
    .Y(_02408_)
  );
  AOI21X1 _08783_ (
    .A(_02546_),
    .B(_02407_),
    .C(_02408_),
    .Y(_01907_)
  );
  AOI22X1 _08784_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_1_ ),
    .Y(_02409_)
  );
  OAI21X1 _08785_ (
    .A(_02170_),
    .B(_02406_),
    .C(_02409_),
    .Y(_01908_)
  );
  AOI22X1 _08786_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_2_ ),
    .Y(_02410_)
  );
  OAI21X1 _08787_ (
    .A(_02172_),
    .B(_02406_),
    .C(_02410_),
    .Y(_01909_)
  );
  AOI22X1 _08788_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_3_ ),
    .Y(_02411_)
  );
  OAI21X1 _08789_ (
    .A(_02177_),
    .B(_02406_),
    .C(_02411_),
    .Y(_01910_)
  );
  AOI22X1 _08790_ (
    .A(_02179_),
    .B(_02405_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_4_ ),
    .Y(_02412_)
  );
  OAI21X1 _08791_ (
    .A(_02559_),
    .B(_02403_),
    .C(_02412_),
    .Y(_01911_)
  );
  AOI22X1 _08792_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_5_ ),
    .Y(_02413_)
  );
  OAI21X1 _08793_ (
    .A(_02184_),
    .B(_02406_),
    .C(_02413_),
    .Y(_01912_)
  );
  AOI22X1 _08794_ (
    .A(_02186_),
    .B(_02405_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_6_ ),
    .Y(_02414_)
  );
  OAI21X1 _08795_ (
    .A(_02562_),
    .B(_02403_),
    .C(_02414_),
    .Y(_01913_)
  );
  AOI22X1 _08796_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_7_ ),
    .Y(_02415_)
  );
  OAI21X1 _08797_ (
    .A(_02191_),
    .B(_02406_),
    .C(_02415_),
    .Y(_01914_)
  );
  AOI22X1 _08798_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_8_ ),
    .Y(_02416_)
  );
  OAI21X1 _08799_ (
    .A(_02193_),
    .B(_02406_),
    .C(_02416_),
    .Y(_01915_)
  );
  AOI22X1 _08800_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_9_ ),
    .Y(_02417_)
  );
  OAI21X1 _08801_ (
    .A(_02198_),
    .B(_02406_),
    .C(_02417_),
    .Y(_01916_)
  );
  AOI22X1 _08802_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_10_ ),
    .Y(_02418_)
  );
  OAI21X1 _08803_ (
    .A(_02200_),
    .B(_02406_),
    .C(_02418_),
    .Y(_01917_)
  );
  AOI22X1 _08804_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_11_ ),
    .Y(_02419_)
  );
  OAI21X1 _08805_ (
    .A(_02205_),
    .B(_02406_),
    .C(_02419_),
    .Y(_01918_)
  );
  AOI22X1 _08806_ (
    .A(_02207_),
    .B(_02405_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_12_ ),
    .Y(_02420_)
  );
  OAI21X1 _08807_ (
    .A(_02739_),
    .B(_02403_),
    .C(_02420_),
    .Y(_01919_)
  );
  AOI22X1 _08808_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_13_ ),
    .Y(_02421_)
  );
  OAI21X1 _08809_ (
    .A(_02212_),
    .B(_02406_),
    .C(_02421_),
    .Y(_01920_)
  );
  AOI22X1 _08810_ (
    .A(_02214_),
    .B(_02405_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_14_ ),
    .Y(_02422_)
  );
  OAI21X1 _08811_ (
    .A(_02767_),
    .B(_02403_),
    .C(_02422_),
    .Y(_01921_)
  );
  AOI22X1 _08812_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02402_),
    .C(_02407_),
    .D( execution_unit_0.register_file_0.r6_15_ ),
    .Y(_02423_)
  );
  OAI21X1 _08813_ (
    .A(_02218_),
    .B(_02406_),
    .C(_02423_),
    .Y(_01922_)
  );
  AND2X1 _08814_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_5_ ),
    .Y(_02424_)
  );
  NAND2X1 _08815_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_5_ ),
    .Y(_02425_)
  );
  NAND2X1 _08816_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02589_),
    .Y(_02426_)
  );
  NOR2X1 _08817_ (
    .A(_02424_),
    .B(_02426_),
    .Y(_02427_)
  );
  OR2X1 _08818_ (
    .A(_02424_),
    .B(_02426_),
    .Y(_02428_)
  );
  AOI21X1 _08819_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02589_),
    .C(_02424_),
    .Y(_02429_)
  );
  OAI22X1 _08820_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .B(_02425_),
    .C(_02428_),
    .D(_02165_),
    .Y(_02430_)
  );
  AOI21X1 _08821_ (
    .A(_02545_),
    .B(_02429_),
    .C(_02430_),
    .Y(_01923_)
  );
  AOI22X1 _08822_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_1_ ),
    .Y(_02431_)
  );
  OAI21X1 _08823_ (
    .A(_02170_),
    .B(_02428_),
    .C(_02431_),
    .Y(_01924_)
  );
  AOI22X1 _08824_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_2_ ),
    .Y(_02432_)
  );
  OAI21X1 _08825_ (
    .A(_02172_),
    .B(_02428_),
    .C(_02432_),
    .Y(_01925_)
  );
  AOI22X1 _08826_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_3_ ),
    .Y(_02433_)
  );
  OAI21X1 _08827_ (
    .A(_02177_),
    .B(_02428_),
    .C(_02433_),
    .Y(_01926_)
  );
  AOI22X1 _08828_ (
    .A(_02179_),
    .B(_02427_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_4_ ),
    .Y(_02434_)
  );
  OAI21X1 _08829_ (
    .A(_02559_),
    .B(_02425_),
    .C(_02434_),
    .Y(_01927_)
  );
  AOI22X1 _08830_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_5_ ),
    .Y(_02435_)
  );
  OAI21X1 _08831_ (
    .A(_02184_),
    .B(_02428_),
    .C(_02435_),
    .Y(_01928_)
  );
  AOI22X1 _08832_ (
    .A(_02186_),
    .B(_02427_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_6_ ),
    .Y(_02436_)
  );
  OAI21X1 _08833_ (
    .A(_02562_),
    .B(_02425_),
    .C(_02436_),
    .Y(_01929_)
  );
  AOI22X1 _08834_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_7_ ),
    .Y(_02437_)
  );
  OAI21X1 _08835_ (
    .A(_02191_),
    .B(_02428_),
    .C(_02437_),
    .Y(_01930_)
  );
  AOI22X1 _08836_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_8_ ),
    .Y(_02438_)
  );
  OAI21X1 _08837_ (
    .A(_02193_),
    .B(_02428_),
    .C(_02438_),
    .Y(_01931_)
  );
  AOI22X1 _08838_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_9_ ),
    .Y(_02439_)
  );
  OAI21X1 _08839_ (
    .A(_02198_),
    .B(_02428_),
    .C(_02439_),
    .Y(_01932_)
  );
  AOI22X1 _08840_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_10_ ),
    .Y(_02440_)
  );
  OAI21X1 _08841_ (
    .A(_02200_),
    .B(_02428_),
    .C(_02440_),
    .Y(_01933_)
  );
  AOI22X1 _08842_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_11_ ),
    .Y(_02441_)
  );
  OAI21X1 _08843_ (
    .A(_02205_),
    .B(_02428_),
    .C(_02441_),
    .Y(_01934_)
  );
  AOI22X1 _08844_ (
    .A(_02207_),
    .B(_02427_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_12_ ),
    .Y(_02442_)
  );
  OAI21X1 _08845_ (
    .A(_02739_),
    .B(_02425_),
    .C(_02442_),
    .Y(_01935_)
  );
  AOI22X1 _08846_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_13_ ),
    .Y(_02443_)
  );
  OAI21X1 _08847_ (
    .A(_02212_),
    .B(_02428_),
    .C(_02443_),
    .Y(_01936_)
  );
  AOI22X1 _08848_ (
    .A(_02214_),
    .B(_02427_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_14_ ),
    .Y(_02444_)
  );
  OAI21X1 _08849_ (
    .A(_02767_),
    .B(_02425_),
    .C(_02444_),
    .Y(_01937_)
  );
  AOI22X1 _08850_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02424_),
    .C(_02429_),
    .D( execution_unit_0.register_file_0.r5_15_ ),
    .Y(_02445_)
  );
  OAI21X1 _08851_ (
    .A(_02218_),
    .B(_02428_),
    .C(_02445_),
    .Y(_01938_)
  );
  AND2X1 _08852_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_4_ ),
    .Y(_02446_)
  );
  NAND2X1 _08853_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_4_ ),
    .Y(_02447_)
  );
  NAND2X1 _08854_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02571_),
    .Y(_02448_)
  );
  NOR2X1 _08855_ (
    .A(_02446_),
    .B(_02448_),
    .Y(_02449_)
  );
  OR2X1 _08856_ (
    .A(_02446_),
    .B(_02448_),
    .Y(_02450_)
  );
  AOI21X1 _08857_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02571_),
    .C(_02446_),
    .Y(_02451_)
  );
  INVX1 _08858_ (
    .A(_02451_),
    .Y(_02452_)
  );
  OAI22X1 _08859_ (
    .A(_02165_),
    .B(_02450_),
    .C(_02452_),
    .D( execution_unit_0.register_file_0.r4_0_ ),
    .Y(_02453_)
  );
  AOI21X1 _08860_ (
    .A(_02551_),
    .B(_02446_),
    .C(_02453_),
    .Y(_01939_)
  );
  AOI22X1 _08861_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_1_ ),
    .Y(_02454_)
  );
  OAI21X1 _08862_ (
    .A(_02170_),
    .B(_02450_),
    .C(_02454_),
    .Y(_01940_)
  );
  AOI22X1 _08863_ (
    .A( execution_unit_0.alu_0.alu_out_2_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_2_ ),
    .Y(_02455_)
  );
  OAI21X1 _08864_ (
    .A(_02172_),
    .B(_02450_),
    .C(_02455_),
    .Y(_01941_)
  );
  AOI22X1 _08865_ (
    .A( execution_unit_0.alu_0.alu_out_3_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_3_ ),
    .Y(_02456_)
  );
  OAI21X1 _08866_ (
    .A(_02177_),
    .B(_02450_),
    .C(_02456_),
    .Y(_01942_)
  );
  AOI22X1 _08867_ (
    .A(_02179_),
    .B(_02449_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_4_ ),
    .Y(_02457_)
  );
  OAI21X1 _08868_ (
    .A(_02559_),
    .B(_02447_),
    .C(_02457_),
    .Y(_01943_)
  );
  AOI22X1 _08869_ (
    .A( execution_unit_0.alu_0.alu_out_5_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_5_ ),
    .Y(_02458_)
  );
  OAI21X1 _08870_ (
    .A(_02184_),
    .B(_02450_),
    .C(_02458_),
    .Y(_01944_)
  );
  AOI22X1 _08871_ (
    .A(_02186_),
    .B(_02449_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_6_ ),
    .Y(_02459_)
  );
  OAI21X1 _08872_ (
    .A(_02562_),
    .B(_02447_),
    .C(_02459_),
    .Y(_01945_)
  );
  AOI22X1 _08873_ (
    .A( execution_unit_0.alu_0.alu_out_7_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_7_ ),
    .Y(_02460_)
  );
  OAI21X1 _08874_ (
    .A(_02191_),
    .B(_02450_),
    .C(_02460_),
    .Y(_01946_)
  );
  AOI22X1 _08875_ (
    .A( execution_unit_0.pc_sw_8_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_8_ ),
    .Y(_02461_)
  );
  OAI21X1 _08876_ (
    .A(_02193_),
    .B(_02450_),
    .C(_02461_),
    .Y(_01947_)
  );
  AOI22X1 _08877_ (
    .A( execution_unit_0.pc_sw_9_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_9_ ),
    .Y(_02462_)
  );
  OAI21X1 _08878_ (
    .A(_02198_),
    .B(_02450_),
    .C(_02462_),
    .Y(_01948_)
  );
  AOI22X1 _08879_ (
    .A( execution_unit_0.pc_sw_10_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_10_ ),
    .Y(_02463_)
  );
  OAI21X1 _08880_ (
    .A(_02200_),
    .B(_02450_),
    .C(_02463_),
    .Y(_01949_)
  );
  AOI22X1 _08881_ (
    .A( execution_unit_0.pc_sw_11_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_11_ ),
    .Y(_02464_)
  );
  OAI21X1 _08882_ (
    .A(_02205_),
    .B(_02450_),
    .C(_02464_),
    .Y(_01950_)
  );
  AOI22X1 _08883_ (
    .A(_02207_),
    .B(_02449_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_12_ ),
    .Y(_02465_)
  );
  OAI21X1 _08884_ (
    .A(_02739_),
    .B(_02447_),
    .C(_02465_),
    .Y(_01951_)
  );
  AOI22X1 _08885_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_13_ ),
    .Y(_02466_)
  );
  OAI21X1 _08886_ (
    .A(_02212_),
    .B(_02450_),
    .C(_02466_),
    .Y(_01952_)
  );
  AOI22X1 _08887_ (
    .A(_02214_),
    .B(_02449_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_14_ ),
    .Y(_02467_)
  );
  OAI21X1 _08888_ (
    .A(_02767_),
    .B(_02447_),
    .C(_02467_),
    .Y(_01953_)
  );
  AOI22X1 _08889_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02446_),
    .C(_02451_),
    .D( execution_unit_0.register_file_0.r4_15_ ),
    .Y(_02468_)
  );
  OAI21X1 _08890_ (
    .A(_02218_),
    .B(_02450_),
    .C(_02468_),
    .Y(_01954_)
  );
  NAND2X1 _08891_ (
    .A( execution_unit_0.reg_dest_wr ),
    .B( execution_unit_0.inst_dest_3_ ),
    .Y(_02469_)
  );
  NAND2X1 _08892_ (
    .A( execution_unit_0.register_file_0.r3_0_ ),
    .B(_02469_),
    .Y(_02470_)
  );
  OAI21X1 _08893_ (
    .A(_02551_),
    .B(_02469_),
    .C(_02470_),
    .Y(_01955_)
  );
  NAND2X1 _08894_ (
    .A( execution_unit_0.register_file_0.r3_1_ ),
    .B(_02469_),
    .Y(_02471_)
  );
  OAI21X1 _08895_ (
    .A(_02554_),
    .B(_02469_),
    .C(_02471_),
    .Y(_01956_)
  );
  NAND2X1 _08896_ (
    .A( execution_unit_0.register_file_0.r3_2_ ),
    .B(_02469_),
    .Y(_02472_)
  );
  OAI21X1 _08897_ (
    .A(_02556_),
    .B(_02469_),
    .C(_02472_),
    .Y(_01957_)
  );
  NAND2X1 _08898_ (
    .A( execution_unit_0.register_file_0.r3_3_ ),
    .B(_02469_),
    .Y(_02473_)
  );
  OAI21X1 _08899_ (
    .A(_02557_),
    .B(_02469_),
    .C(_02473_),
    .Y(_01958_)
  );
  NAND2X1 _08900_ (
    .A( execution_unit_0.register_file_0.r3_4_ ),
    .B(_02469_),
    .Y(_02474_)
  );
  OAI21X1 _08901_ (
    .A(_02559_),
    .B(_02469_),
    .C(_02474_),
    .Y(_01959_)
  );
  NAND2X1 _08902_ (
    .A( execution_unit_0.register_file_0.r3_5_ ),
    .B(_02469_),
    .Y(_02475_)
  );
  OAI21X1 _08903_ (
    .A(_02561_),
    .B(_02469_),
    .C(_02475_),
    .Y(_01960_)
  );
  NAND2X1 _08904_ (
    .A( execution_unit_0.register_file_0.r3_6_ ),
    .B(_02469_),
    .Y(_02476_)
  );
  OAI21X1 _08905_ (
    .A(_02562_),
    .B(_02469_),
    .C(_02476_),
    .Y(_01961_)
  );
  NAND2X1 _08906_ (
    .A( execution_unit_0.register_file_0.r3_7_ ),
    .B(_02469_),
    .Y(_02477_)
  );
  OAI21X1 _08907_ (
    .A(_02563_),
    .B(_02469_),
    .C(_02477_),
    .Y(_01962_)
  );
  NAND2X1 _08908_ (
    .A( execution_unit_0.register_file_0.r3_8_ ),
    .B(_02469_),
    .Y(_02478_)
  );
  OAI21X1 _08909_ (
    .A(_02678_),
    .B(_02469_),
    .C(_02478_),
    .Y(_01963_)
  );
  NAND2X1 _08910_ (
    .A( execution_unit_0.register_file_0.r3_9_ ),
    .B(_02469_),
    .Y(_02479_)
  );
  OAI21X1 _08911_ (
    .A(_02694_),
    .B(_02469_),
    .C(_02479_),
    .Y(_01964_)
  );
  NAND2X1 _08912_ (
    .A( execution_unit_0.register_file_0.r3_10_ ),
    .B(_02469_),
    .Y(_02480_)
  );
  OAI21X1 _08913_ (
    .A(_02709_),
    .B(_02469_),
    .C(_02480_),
    .Y(_01965_)
  );
  NAND2X1 _08914_ (
    .A( execution_unit_0.register_file_0.r3_11_ ),
    .B(_02469_),
    .Y(_02481_)
  );
  OAI21X1 _08915_ (
    .A(_02725_),
    .B(_02469_),
    .C(_02481_),
    .Y(_01966_)
  );
  NAND2X1 _08916_ (
    .A( execution_unit_0.register_file_0.r3_12_ ),
    .B(_02469_),
    .Y(_02482_)
  );
  OAI21X1 _08917_ (
    .A(_02739_),
    .B(_02469_),
    .C(_02482_),
    .Y(_01967_)
  );
  NAND2X1 _08918_ (
    .A( execution_unit_0.register_file_0.r3_13_ ),
    .B(_02469_),
    .Y(_02483_)
  );
  OAI21X1 _08919_ (
    .A(_02753_),
    .B(_02469_),
    .C(_02483_),
    .Y(_01968_)
  );
  NAND2X1 _08920_ (
    .A( execution_unit_0.register_file_0.r3_14_ ),
    .B(_02469_),
    .Y(_02484_)
  );
  OAI21X1 _08921_ (
    .A(_02767_),
    .B(_02469_),
    .C(_02484_),
    .Y(_01969_)
  );
  NAND2X1 _08922_ (
    .A( execution_unit_0.register_file_0.r3_15_ ),
    .B(_02469_),
    .Y(_02485_)
  );
  OAI21X1 _08923_ (
    .A(_02782_),
    .B(_02469_),
    .C(_02485_),
    .Y(_01970_)
  );
  NOR2X1 _08924_ (
    .A(_02551_),
    .B(_02795_),
    .Y(_02486_)
  );
  AOI22X1 _08925_ (
    .A( execution_unit_0.alu_0.status_0_ ),
    .B(_02146_),
    .C(_02486_),
    .D(_02540_),
    .Y(_02487_)
  );
  NAND3X1 _08926_ (
    .A(_02540_),
    .B( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .C( execution_unit_0.alu_0.alu_stat_0_ ),
    .Y(_02488_)
  );
  OAI21X1 _08927_ (
    .A( execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .B(_02487_),
    .C(_02488_),
    .Y(_01971_)
  );
  AND2X1 _08928_ (
    .A(_02539_),
    .B(_02170_),
    .Y(_02489_)
  );
  AND2X1 _08929_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.reg_dest_wr ),
    .Y(_02490_)
  );
  NAND2X1 _08930_ (
    .A( execution_unit_0.inst_dest_1_ ),
    .B( execution_unit_0.reg_dest_wr ),
    .Y(_02491_)
  );
  AOI21X1 _08931_ (
    .A( execution_unit_0.reg_incr ),
    .B(_02566_),
    .C( execution_unit_0.reg_sp_wr ),
    .Y(_02492_)
  );
  NOR2X1 _08932_ (
    .A(_02490_),
    .B(_02492_),
    .Y(_02493_)
  );
  OAI21X1 _08933_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_1_ ),
    .C(_02493_),
    .Y(_02494_)
  );
  AND2X1 _08934_ (
    .A(_02491_),
    .B(_02492_),
    .Y(_02495_)
  );
  AOI22X1 _08935_ (
    .A( execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_1_ ),
    .Y(_02496_)
  );
  OAI21X1 _08936_ (
    .A(_02489_),
    .B(_02494_),
    .C(_02496_),
    .Y(_01972_)
  );
  OAI21X1 _08937_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_2_ ),
    .C(_02493_),
    .Y(_02497_)
  );
  AOI21X1 _08938_ (
    .A(_02539_),
    .B(_02172_),
    .C(_02497_),
    .Y(_02498_)
  );
  AOI21X1 _08939_ (
    .A( execution_unit_0.register_file_0.r1_2_ ),
    .B(_02495_),
    .C(_02498_),
    .Y(_02499_)
  );
  OAI21X1 _08940_ (
    .A(_02556_),
    .B(_02491_),
    .C(_02499_),
    .Y(_01973_)
  );
  OAI21X1 _08941_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_3_ ),
    .C(_02493_),
    .Y(_02500_)
  );
  AOI21X1 _08942_ (
    .A(_02539_),
    .B(_02177_),
    .C(_02500_),
    .Y(_02501_)
  );
  AOI21X1 _08943_ (
    .A( execution_unit_0.register_file_0.r1_3_ ),
    .B(_02495_),
    .C(_02501_),
    .Y(_02502_)
  );
  OAI21X1 _08944_ (
    .A(_02557_),
    .B(_02491_),
    .C(_02502_),
    .Y(_01974_)
  );
  NOR2X1 _08945_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02179_),
    .Y(_02503_)
  );
  OAI21X1 _08946_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_4_ ),
    .C(_02493_),
    .Y(_02504_)
  );
  AOI22X1 _08947_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_4_ ),
    .Y(_02505_)
  );
  OAI21X1 _08948_ (
    .A(_02503_),
    .B(_02504_),
    .C(_02505_),
    .Y(_01975_)
  );
  OAI21X1 _08949_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_5_ ),
    .C(_02493_),
    .Y(_02506_)
  );
  AOI21X1 _08950_ (
    .A(_02539_),
    .B(_02184_),
    .C(_02506_),
    .Y(_02507_)
  );
  AOI21X1 _08951_ (
    .A( execution_unit_0.register_file_0.r1_5_ ),
    .B(_02495_),
    .C(_02507_),
    .Y(_02508_)
  );
  OAI21X1 _08952_ (
    .A(_02561_),
    .B(_02491_),
    .C(_02508_),
    .Y(_01976_)
  );
  NOR2X1 _08953_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02186_),
    .Y(_02509_)
  );
  OAI21X1 _08954_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_6_ ),
    .C(_02493_),
    .Y(_02510_)
  );
  AOI22X1 _08955_ (
    .A( execution_unit_0.alu_0.alu_out_6_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_6_ ),
    .Y(_02511_)
  );
  OAI21X1 _08956_ (
    .A(_02509_),
    .B(_02510_),
    .C(_02511_),
    .Y(_01977_)
  );
  OAI21X1 _08957_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_7_ ),
    .C(_02493_),
    .Y(_02512_)
  );
  AOI21X1 _08958_ (
    .A(_02539_),
    .B(_02191_),
    .C(_02512_),
    .Y(_02513_)
  );
  AOI21X1 _08959_ (
    .A( execution_unit_0.register_file_0.r1_7_ ),
    .B(_02495_),
    .C(_02513_),
    .Y(_02514_)
  );
  OAI21X1 _08960_ (
    .A(_02563_),
    .B(_02491_),
    .C(_02514_),
    .Y(_01978_)
  );
  OAI21X1 _08961_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_8_ ),
    .C(_02493_),
    .Y(_02515_)
  );
  AOI21X1 _08962_ (
    .A(_02539_),
    .B(_02193_),
    .C(_02515_),
    .Y(_02516_)
  );
  AOI21X1 _08963_ (
    .A( execution_unit_0.register_file_0.r1_8_ ),
    .B(_02495_),
    .C(_02516_),
    .Y(_02517_)
  );
  OAI21X1 _08964_ (
    .A(_02678_),
    .B(_02491_),
    .C(_02517_),
    .Y(_01979_)
  );
  OAI21X1 _08965_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_9_ ),
    .C(_02493_),
    .Y(_02518_)
  );
  AOI21X1 _08966_ (
    .A(_02539_),
    .B(_02198_),
    .C(_02518_),
    .Y(_02519_)
  );
  AOI21X1 _08967_ (
    .A( execution_unit_0.register_file_0.r1_9_ ),
    .B(_02495_),
    .C(_02519_),
    .Y(_02520_)
  );
  OAI21X1 _08968_ (
    .A(_02694_),
    .B(_02491_),
    .C(_02520_),
    .Y(_01980_)
  );
  OAI21X1 _08969_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_10_ ),
    .C(_02493_),
    .Y(_02521_)
  );
  AOI21X1 _08970_ (
    .A(_02539_),
    .B(_02200_),
    .C(_02521_),
    .Y(_02522_)
  );
  AOI21X1 _08971_ (
    .A( execution_unit_0.register_file_0.r1_10_ ),
    .B(_02495_),
    .C(_02522_),
    .Y(_02523_)
  );
  OAI21X1 _08972_ (
    .A(_02709_),
    .B(_02491_),
    .C(_02523_),
    .Y(_01981_)
  );
  OAI21X1 _08973_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_11_ ),
    .C(_02493_),
    .Y(_02524_)
  );
  AOI21X1 _08974_ (
    .A(_02539_),
    .B(_02205_),
    .C(_02524_),
    .Y(_02525_)
  );
  AOI21X1 _08975_ (
    .A( execution_unit_0.register_file_0.r1_11_ ),
    .B(_02495_),
    .C(_02525_),
    .Y(_02526_)
  );
  OAI21X1 _08976_ (
    .A(_02725_),
    .B(_02491_),
    .C(_02526_),
    .Y(_01982_)
  );
  NOR2X1 _08977_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02207_),
    .Y(_02527_)
  );
  OAI21X1 _08978_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_12_ ),
    .C(_02493_),
    .Y(_02528_)
  );
  AOI22X1 _08979_ (
    .A( execution_unit_0.pc_sw_12_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_12_ ),
    .Y(_02529_)
  );
  OAI21X1 _08980_ (
    .A(_02527_),
    .B(_02528_),
    .C(_02529_),
    .Y(_01983_)
  );
  AOI21X1 _08981_ (
    .A(_02210_),
    .B(_02211_),
    .C( execution_unit_0.reg_sp_wr ),
    .Y(_02530_)
  );
  OAI21X1 _08982_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_13_ ),
    .C(_02493_),
    .Y(_02531_)
  );
  AOI22X1 _08983_ (
    .A( execution_unit_0.pc_sw_13_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_13_ ),
    .Y(_02532_)
  );
  OAI21X1 _08984_ (
    .A(_02530_),
    .B(_02531_),
    .C(_02532_),
    .Y(_01984_)
  );
  NOR2X1 _08985_ (
    .A( execution_unit_0.reg_sp_wr ),
    .B(_02214_),
    .Y(_02533_)
  );
  OAI21X1 _08986_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .C(_02493_),
    .Y(_02534_)
  );
  AOI22X1 _08987_ (
    .A( execution_unit_0.pc_sw_14_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_14_ ),
    .Y(_02535_)
  );
  OAI21X1 _08988_ (
    .A(_02533_),
    .B(_02534_),
    .C(_02535_),
    .Y(_01985_)
  );
  AOI21X1 _08989_ (
    .A(_02216_),
    .B(_02217_),
    .C( execution_unit_0.reg_sp_wr ),
    .Y(_02536_)
  );
  OAI21X1 _08990_ (
    .A(_02539_),
    .B( dbg_0.UNUSED_eu_mab_15_ ),
    .C(_02493_),
    .Y(_02537_)
  );
  AOI22X1 _08991_ (
    .A( execution_unit_0.pc_sw_15_ ),
    .B(_02490_),
    .C(_02495_),
    .D( execution_unit_0.register_file_0.r1_15_ ),
    .Y(_02538_)
  );
  OAI21X1 _08992_ (
    .A(_02536_),
    .B(_02537_),
    .C(_02538_),
    .Y(_01986_)
  );
  DFFSR _08993_ (
    .CLK(dco_clk),
    .D(_01757_),
    .Q( execution_unit_0.alu_0.status_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _08994_ (
    .CLK(dco_clk),
    .D(_01758_),
    .Q( execution_unit_0.alu_0.status_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _08995_ (
    .CLK(dco_clk),
    .D(_01759_),
    .Q( execution_unit_0.gie ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _08996_ (
    .CLK(dco_clk),
    .D(_01760_),
    .Q( clock_module_0.oscoff ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _08997_ (
    .CLK(dco_clk),
    .D(_01761_),
    .Q( clock_module_0.scg1 ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _08998_ (
    .CLK(dco_clk),
    .D(_01762_),
    .Q( execution_unit_0.alu_0.status_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _08999_ (
    .CLK(dco_clk),
    .D(_01763_),
    .Q( execution_unit_0.register_file_0.r15_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09000_ (
    .CLK(dco_clk),
    .D(_01764_),
    .Q( execution_unit_0.register_file_0.r15_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09001_ (
    .CLK(dco_clk),
    .D(_01765_),
    .Q( execution_unit_0.register_file_0.r15_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09002_ (
    .CLK(dco_clk),
    .D(_01766_),
    .Q( execution_unit_0.register_file_0.r15_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09003_ (
    .CLK(dco_clk),
    .D(_01767_),
    .Q( execution_unit_0.register_file_0.r15_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09004_ (
    .CLK(dco_clk),
    .D(_01768_),
    .Q( execution_unit_0.register_file_0.r15_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09005_ (
    .CLK(dco_clk),
    .D(_01769_),
    .Q( execution_unit_0.register_file_0.r15_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09006_ (
    .CLK(dco_clk),
    .D(_01770_),
    .Q( execution_unit_0.register_file_0.r15_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09007_ (
    .CLK(dco_clk),
    .D(_01771_),
    .Q( execution_unit_0.register_file_0.r15_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09008_ (
    .CLK(dco_clk),
    .D(_01772_),
    .Q( execution_unit_0.register_file_0.r15_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09009_ (
    .CLK(dco_clk),
    .D(_01773_),
    .Q( execution_unit_0.register_file_0.r15_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09010_ (
    .CLK(dco_clk),
    .D(_01774_),
    .Q( execution_unit_0.register_file_0.r15_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09011_ (
    .CLK(dco_clk),
    .D(_01775_),
    .Q( execution_unit_0.register_file_0.r15_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09012_ (
    .CLK(dco_clk),
    .D(_01776_),
    .Q( execution_unit_0.register_file_0.r15_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09013_ (
    .CLK(dco_clk),
    .D(_01777_),
    .Q( execution_unit_0.register_file_0.r15_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09014_ (
    .CLK(dco_clk),
    .D(_01778_),
    .Q( execution_unit_0.register_file_0.r15_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09015_ (
    .CLK(dco_clk),
    .D(_01779_),
    .Q( execution_unit_0.register_file_0.r14_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09016_ (
    .CLK(dco_clk),
    .D(_01780_),
    .Q( execution_unit_0.register_file_0.r14_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09017_ (
    .CLK(dco_clk),
    .D(_01781_),
    .Q( execution_unit_0.register_file_0.r14_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09018_ (
    .CLK(dco_clk),
    .D(_01782_),
    .Q( execution_unit_0.register_file_0.r14_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09019_ (
    .CLK(dco_clk),
    .D(_01783_),
    .Q( execution_unit_0.register_file_0.r14_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09020_ (
    .CLK(dco_clk),
    .D(_01784_),
    .Q( execution_unit_0.register_file_0.r14_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09021_ (
    .CLK(dco_clk),
    .D(_01785_),
    .Q( execution_unit_0.register_file_0.r14_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09022_ (
    .CLK(dco_clk),
    .D(_01786_),
    .Q( execution_unit_0.register_file_0.r14_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09023_ (
    .CLK(dco_clk),
    .D(_01787_),
    .Q( execution_unit_0.register_file_0.r14_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09024_ (
    .CLK(dco_clk),
    .D(_01788_),
    .Q( execution_unit_0.register_file_0.r14_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09025_ (
    .CLK(dco_clk),
    .D(_01789_),
    .Q( execution_unit_0.register_file_0.r14_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09026_ (
    .CLK(dco_clk),
    .D(_01790_),
    .Q( execution_unit_0.register_file_0.r14_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09027_ (
    .CLK(dco_clk),
    .D(_01791_),
    .Q( execution_unit_0.register_file_0.r14_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09028_ (
    .CLK(dco_clk),
    .D(_01792_),
    .Q( execution_unit_0.register_file_0.r14_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09029_ (
    .CLK(dco_clk),
    .D(_01793_),
    .Q( execution_unit_0.register_file_0.r14_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09030_ (
    .CLK(dco_clk),
    .D(_01794_),
    .Q( execution_unit_0.register_file_0.r14_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09031_ (
    .CLK(dco_clk),
    .D(_01795_),
    .Q( execution_unit_0.register_file_0.r13_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09032_ (
    .CLK(dco_clk),
    .D(_01796_),
    .Q( execution_unit_0.register_file_0.r13_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09033_ (
    .CLK(dco_clk),
    .D(_01797_),
    .Q( execution_unit_0.register_file_0.r13_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09034_ (
    .CLK(dco_clk),
    .D(_01798_),
    .Q( execution_unit_0.register_file_0.r13_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09035_ (
    .CLK(dco_clk),
    .D(_01799_),
    .Q( execution_unit_0.register_file_0.r13_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09036_ (
    .CLK(dco_clk),
    .D(_01800_),
    .Q( execution_unit_0.register_file_0.r13_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09037_ (
    .CLK(dco_clk),
    .D(_01801_),
    .Q( execution_unit_0.register_file_0.r13_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09038_ (
    .CLK(dco_clk),
    .D(_01802_),
    .Q( execution_unit_0.register_file_0.r13_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09039_ (
    .CLK(dco_clk),
    .D(_01803_),
    .Q( execution_unit_0.register_file_0.r13_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09040_ (
    .CLK(dco_clk),
    .D(_01804_),
    .Q( execution_unit_0.register_file_0.r13_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09041_ (
    .CLK(dco_clk),
    .D(_01805_),
    .Q( execution_unit_0.register_file_0.r13_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09042_ (
    .CLK(dco_clk),
    .D(_01806_),
    .Q( execution_unit_0.register_file_0.r13_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09043_ (
    .CLK(dco_clk),
    .D(_01807_),
    .Q( execution_unit_0.register_file_0.r13_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09044_ (
    .CLK(dco_clk),
    .D(_01808_),
    .Q( execution_unit_0.register_file_0.r13_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09045_ (
    .CLK(dco_clk),
    .D(_01809_),
    .Q( execution_unit_0.register_file_0.r13_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09046_ (
    .CLK(dco_clk),
    .D(_01810_),
    .Q( execution_unit_0.register_file_0.r13_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09047_ (
    .CLK(dco_clk),
    .D(_01811_),
    .Q( execution_unit_0.register_file_0.r12_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09048_ (
    .CLK(dco_clk),
    .D(_01812_),
    .Q( execution_unit_0.register_file_0.r12_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09049_ (
    .CLK(dco_clk),
    .D(_01813_),
    .Q( execution_unit_0.register_file_0.r12_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09050_ (
    .CLK(dco_clk),
    .D(_01814_),
    .Q( execution_unit_0.register_file_0.r12_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09051_ (
    .CLK(dco_clk),
    .D(_01815_),
    .Q( execution_unit_0.register_file_0.r12_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09052_ (
    .CLK(dco_clk),
    .D(_01816_),
    .Q( execution_unit_0.register_file_0.r12_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09053_ (
    .CLK(dco_clk),
    .D(_01817_),
    .Q( execution_unit_0.register_file_0.r12_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09054_ (
    .CLK(dco_clk),
    .D(_01818_),
    .Q( execution_unit_0.register_file_0.r12_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09055_ (
    .CLK(dco_clk),
    .D(_01819_),
    .Q( execution_unit_0.register_file_0.r12_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09056_ (
    .CLK(dco_clk),
    .D(_01820_),
    .Q( execution_unit_0.register_file_0.r12_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09057_ (
    .CLK(dco_clk),
    .D(_01821_),
    .Q( execution_unit_0.register_file_0.r12_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09058_ (
    .CLK(dco_clk),
    .D(_01822_),
    .Q( execution_unit_0.register_file_0.r12_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09059_ (
    .CLK(dco_clk),
    .D(_01823_),
    .Q( execution_unit_0.register_file_0.r12_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09060_ (
    .CLK(dco_clk),
    .D(_01824_),
    .Q( execution_unit_0.register_file_0.r12_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09061_ (
    .CLK(dco_clk),
    .D(_01825_),
    .Q( execution_unit_0.register_file_0.r12_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09062_ (
    .CLK(dco_clk),
    .D(_01826_),
    .Q( execution_unit_0.register_file_0.r12_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09063_ (
    .CLK(dco_clk),
    .D(_01827_),
    .Q( execution_unit_0.register_file_0.r11_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09064_ (
    .CLK(dco_clk),
    .D(_01828_),
    .Q( execution_unit_0.register_file_0.r11_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09065_ (
    .CLK(dco_clk),
    .D(_01829_),
    .Q( execution_unit_0.register_file_0.r11_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09066_ (
    .CLK(dco_clk),
    .D(_01830_),
    .Q( execution_unit_0.register_file_0.r11_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09067_ (
    .CLK(dco_clk),
    .D(_01831_),
    .Q( execution_unit_0.register_file_0.r11_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09068_ (
    .CLK(dco_clk),
    .D(_01832_),
    .Q( execution_unit_0.register_file_0.r11_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09069_ (
    .CLK(dco_clk),
    .D(_01833_),
    .Q( execution_unit_0.register_file_0.r11_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09070_ (
    .CLK(dco_clk),
    .D(_01834_),
    .Q( execution_unit_0.register_file_0.r11_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09071_ (
    .CLK(dco_clk),
    .D(_01835_),
    .Q( execution_unit_0.register_file_0.r11_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09072_ (
    .CLK(dco_clk),
    .D(_01836_),
    .Q( execution_unit_0.register_file_0.r11_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09073_ (
    .CLK(dco_clk),
    .D(_01837_),
    .Q( execution_unit_0.register_file_0.r11_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09074_ (
    .CLK(dco_clk),
    .D(_01838_),
    .Q( execution_unit_0.register_file_0.r11_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09075_ (
    .CLK(dco_clk),
    .D(_01839_),
    .Q( execution_unit_0.register_file_0.r11_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09076_ (
    .CLK(dco_clk),
    .D(_01840_),
    .Q( execution_unit_0.register_file_0.r11_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09077_ (
    .CLK(dco_clk),
    .D(_01841_),
    .Q( execution_unit_0.register_file_0.r11_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09078_ (
    .CLK(dco_clk),
    .D(_01842_),
    .Q( execution_unit_0.register_file_0.r11_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09079_ (
    .CLK(dco_clk),
    .D(_01843_),
    .Q( execution_unit_0.register_file_0.r10_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09080_ (
    .CLK(dco_clk),
    .D(_01844_),
    .Q( execution_unit_0.register_file_0.r10_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09081_ (
    .CLK(dco_clk),
    .D(_01845_),
    .Q( execution_unit_0.register_file_0.r10_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09082_ (
    .CLK(dco_clk),
    .D(_01846_),
    .Q( execution_unit_0.register_file_0.r10_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09083_ (
    .CLK(dco_clk),
    .D(_01847_),
    .Q( execution_unit_0.register_file_0.r10_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09084_ (
    .CLK(dco_clk),
    .D(_01848_),
    .Q( execution_unit_0.register_file_0.r10_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09085_ (
    .CLK(dco_clk),
    .D(_01849_),
    .Q( execution_unit_0.register_file_0.r10_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09086_ (
    .CLK(dco_clk),
    .D(_01850_),
    .Q( execution_unit_0.register_file_0.r10_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09087_ (
    .CLK(dco_clk),
    .D(_01851_),
    .Q( execution_unit_0.register_file_0.r10_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09088_ (
    .CLK(dco_clk),
    .D(_01852_),
    .Q( execution_unit_0.register_file_0.r10_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09089_ (
    .CLK(dco_clk),
    .D(_01853_),
    .Q( execution_unit_0.register_file_0.r10_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09090_ (
    .CLK(dco_clk),
    .D(_01854_),
    .Q( execution_unit_0.register_file_0.r10_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09091_ (
    .CLK(dco_clk),
    .D(_01855_),
    .Q( execution_unit_0.register_file_0.r10_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09092_ (
    .CLK(dco_clk),
    .D(_01856_),
    .Q( execution_unit_0.register_file_0.r10_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09093_ (
    .CLK(dco_clk),
    .D(_01857_),
    .Q( execution_unit_0.register_file_0.r10_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09094_ (
    .CLK(dco_clk),
    .D(_01858_),
    .Q( execution_unit_0.register_file_0.r10_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09095_ (
    .CLK(dco_clk),
    .D(_01859_),
    .Q( execution_unit_0.register_file_0.r9_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09096_ (
    .CLK(dco_clk),
    .D(_01860_),
    .Q( execution_unit_0.register_file_0.r9_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09097_ (
    .CLK(dco_clk),
    .D(_01861_),
    .Q( execution_unit_0.register_file_0.r9_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09098_ (
    .CLK(dco_clk),
    .D(_01862_),
    .Q( execution_unit_0.register_file_0.r9_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09099_ (
    .CLK(dco_clk),
    .D(_01863_),
    .Q( execution_unit_0.register_file_0.r9_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09100_ (
    .CLK(dco_clk),
    .D(_01864_),
    .Q( execution_unit_0.register_file_0.r9_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09101_ (
    .CLK(dco_clk),
    .D(_01865_),
    .Q( execution_unit_0.register_file_0.r9_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09102_ (
    .CLK(dco_clk),
    .D(_01866_),
    .Q( execution_unit_0.register_file_0.r9_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09103_ (
    .CLK(dco_clk),
    .D(_01867_),
    .Q( execution_unit_0.register_file_0.r9_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09104_ (
    .CLK(dco_clk),
    .D(_01868_),
    .Q( execution_unit_0.register_file_0.r9_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09105_ (
    .CLK(dco_clk),
    .D(_01869_),
    .Q( execution_unit_0.register_file_0.r9_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09106_ (
    .CLK(dco_clk),
    .D(_01870_),
    .Q( execution_unit_0.register_file_0.r9_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09107_ (
    .CLK(dco_clk),
    .D(_01871_),
    .Q( execution_unit_0.register_file_0.r9_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09108_ (
    .CLK(dco_clk),
    .D(_01872_),
    .Q( execution_unit_0.register_file_0.r9_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09109_ (
    .CLK(dco_clk),
    .D(_01873_),
    .Q( execution_unit_0.register_file_0.r9_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09110_ (
    .CLK(dco_clk),
    .D(_01874_),
    .Q( execution_unit_0.register_file_0.r9_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09111_ (
    .CLK(dco_clk),
    .D(_01875_),
    .Q( execution_unit_0.register_file_0.r8_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09112_ (
    .CLK(dco_clk),
    .D(_01876_),
    .Q( execution_unit_0.register_file_0.r8_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09113_ (
    .CLK(dco_clk),
    .D(_01877_),
    .Q( execution_unit_0.register_file_0.r8_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09114_ (
    .CLK(dco_clk),
    .D(_01878_),
    .Q( execution_unit_0.register_file_0.r8_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09115_ (
    .CLK(dco_clk),
    .D(_01879_),
    .Q( execution_unit_0.register_file_0.r8_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09116_ (
    .CLK(dco_clk),
    .D(_01880_),
    .Q( execution_unit_0.register_file_0.r8_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09117_ (
    .CLK(dco_clk),
    .D(_01881_),
    .Q( execution_unit_0.register_file_0.r8_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09118_ (
    .CLK(dco_clk),
    .D(_01882_),
    .Q( execution_unit_0.register_file_0.r8_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09119_ (
    .CLK(dco_clk),
    .D(_01883_),
    .Q( execution_unit_0.register_file_0.r8_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09120_ (
    .CLK(dco_clk),
    .D(_01884_),
    .Q( execution_unit_0.register_file_0.r8_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09121_ (
    .CLK(dco_clk),
    .D(_01885_),
    .Q( execution_unit_0.register_file_0.r8_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09122_ (
    .CLK(dco_clk),
    .D(_01886_),
    .Q( execution_unit_0.register_file_0.r8_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09123_ (
    .CLK(dco_clk),
    .D(_01887_),
    .Q( execution_unit_0.register_file_0.r8_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09124_ (
    .CLK(dco_clk),
    .D(_01888_),
    .Q( execution_unit_0.register_file_0.r8_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09125_ (
    .CLK(dco_clk),
    .D(_01889_),
    .Q( execution_unit_0.register_file_0.r8_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09126_ (
    .CLK(dco_clk),
    .D(_01890_),
    .Q( execution_unit_0.register_file_0.r8_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09127_ (
    .CLK(dco_clk),
    .D(_01891_),
    .Q( execution_unit_0.register_file_0.r7_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09128_ (
    .CLK(dco_clk),
    .D(_01892_),
    .Q( execution_unit_0.register_file_0.r7_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09129_ (
    .CLK(dco_clk),
    .D(_01893_),
    .Q( execution_unit_0.register_file_0.r7_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09130_ (
    .CLK(dco_clk),
    .D(_01894_),
    .Q( execution_unit_0.register_file_0.r7_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09131_ (
    .CLK(dco_clk),
    .D(_01895_),
    .Q( execution_unit_0.register_file_0.r7_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09132_ (
    .CLK(dco_clk),
    .D(_01896_),
    .Q( execution_unit_0.register_file_0.r7_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09133_ (
    .CLK(dco_clk),
    .D(_01897_),
    .Q( execution_unit_0.register_file_0.r7_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09134_ (
    .CLK(dco_clk),
    .D(_01898_),
    .Q( execution_unit_0.register_file_0.r7_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09135_ (
    .CLK(dco_clk),
    .D(_01899_),
    .Q( execution_unit_0.register_file_0.r7_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09136_ (
    .CLK(dco_clk),
    .D(_01900_),
    .Q( execution_unit_0.register_file_0.r7_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09137_ (
    .CLK(dco_clk),
    .D(_01901_),
    .Q( execution_unit_0.register_file_0.r7_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09138_ (
    .CLK(dco_clk),
    .D(_01902_),
    .Q( execution_unit_0.register_file_0.r7_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09139_ (
    .CLK(dco_clk),
    .D(_01903_),
    .Q( execution_unit_0.register_file_0.r7_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09140_ (
    .CLK(dco_clk),
    .D(_01904_),
    .Q( execution_unit_0.register_file_0.r7_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09141_ (
    .CLK(dco_clk),
    .D(_01905_),
    .Q( execution_unit_0.register_file_0.r7_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09142_ (
    .CLK(dco_clk),
    .D(_01906_),
    .Q( execution_unit_0.register_file_0.r7_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09143_ (
    .CLK(dco_clk),
    .D(_01907_),
    .Q( execution_unit_0.register_file_0.r6_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09144_ (
    .CLK(dco_clk),
    .D(_01908_),
    .Q( execution_unit_0.register_file_0.r6_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09145_ (
    .CLK(dco_clk),
    .D(_01909_),
    .Q( execution_unit_0.register_file_0.r6_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09146_ (
    .CLK(dco_clk),
    .D(_01910_),
    .Q( execution_unit_0.register_file_0.r6_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09147_ (
    .CLK(dco_clk),
    .D(_01911_),
    .Q( execution_unit_0.register_file_0.r6_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09148_ (
    .CLK(dco_clk),
    .D(_01912_),
    .Q( execution_unit_0.register_file_0.r6_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09149_ (
    .CLK(dco_clk),
    .D(_01913_),
    .Q( execution_unit_0.register_file_0.r6_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09150_ (
    .CLK(dco_clk),
    .D(_01914_),
    .Q( execution_unit_0.register_file_0.r6_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09151_ (
    .CLK(dco_clk),
    .D(_01915_),
    .Q( execution_unit_0.register_file_0.r6_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09152_ (
    .CLK(dco_clk),
    .D(_01916_),
    .Q( execution_unit_0.register_file_0.r6_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09153_ (
    .CLK(dco_clk),
    .D(_01917_),
    .Q( execution_unit_0.register_file_0.r6_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09154_ (
    .CLK(dco_clk),
    .D(_01918_),
    .Q( execution_unit_0.register_file_0.r6_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09155_ (
    .CLK(dco_clk),
    .D(_01919_),
    .Q( execution_unit_0.register_file_0.r6_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09156_ (
    .CLK(dco_clk),
    .D(_01920_),
    .Q( execution_unit_0.register_file_0.r6_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09157_ (
    .CLK(dco_clk),
    .D(_01921_),
    .Q( execution_unit_0.register_file_0.r6_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09158_ (
    .CLK(dco_clk),
    .D(_01922_),
    .Q( execution_unit_0.register_file_0.r6_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09159_ (
    .CLK(dco_clk),
    .D(_01923_),
    .Q( execution_unit_0.register_file_0.r5_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09160_ (
    .CLK(dco_clk),
    .D(_01924_),
    .Q( execution_unit_0.register_file_0.r5_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09161_ (
    .CLK(dco_clk),
    .D(_01925_),
    .Q( execution_unit_0.register_file_0.r5_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09162_ (
    .CLK(dco_clk),
    .D(_01926_),
    .Q( execution_unit_0.register_file_0.r5_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09163_ (
    .CLK(dco_clk),
    .D(_01927_),
    .Q( execution_unit_0.register_file_0.r5_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09164_ (
    .CLK(dco_clk),
    .D(_01928_),
    .Q( execution_unit_0.register_file_0.r5_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09165_ (
    .CLK(dco_clk),
    .D(_01929_),
    .Q( execution_unit_0.register_file_0.r5_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09166_ (
    .CLK(dco_clk),
    .D(_01930_),
    .Q( execution_unit_0.register_file_0.r5_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09167_ (
    .CLK(dco_clk),
    .D(_01931_),
    .Q( execution_unit_0.register_file_0.r5_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09168_ (
    .CLK(dco_clk),
    .D(_01932_),
    .Q( execution_unit_0.register_file_0.r5_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09169_ (
    .CLK(dco_clk),
    .D(_01933_),
    .Q( execution_unit_0.register_file_0.r5_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09170_ (
    .CLK(dco_clk),
    .D(_01934_),
    .Q( execution_unit_0.register_file_0.r5_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09171_ (
    .CLK(dco_clk),
    .D(_01935_),
    .Q( execution_unit_0.register_file_0.r5_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09172_ (
    .CLK(dco_clk),
    .D(_01936_),
    .Q( execution_unit_0.register_file_0.r5_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09173_ (
    .CLK(dco_clk),
    .D(_01937_),
    .Q( execution_unit_0.register_file_0.r5_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09174_ (
    .CLK(dco_clk),
    .D(_01938_),
    .Q( execution_unit_0.register_file_0.r5_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09175_ (
    .CLK(dco_clk),
    .D(_01939_),
    .Q( execution_unit_0.register_file_0.r4_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09176_ (
    .CLK(dco_clk),
    .D(_01940_),
    .Q( execution_unit_0.register_file_0.r4_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09177_ (
    .CLK(dco_clk),
    .D(_01941_),
    .Q( execution_unit_0.register_file_0.r4_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09178_ (
    .CLK(dco_clk),
    .D(_01942_),
    .Q( execution_unit_0.register_file_0.r4_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09179_ (
    .CLK(dco_clk),
    .D(_01943_),
    .Q( execution_unit_0.register_file_0.r4_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09180_ (
    .CLK(dco_clk),
    .D(_01944_),
    .Q( execution_unit_0.register_file_0.r4_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09181_ (
    .CLK(dco_clk),
    .D(_01945_),
    .Q( execution_unit_0.register_file_0.r4_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09182_ (
    .CLK(dco_clk),
    .D(_01946_),
    .Q( execution_unit_0.register_file_0.r4_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09183_ (
    .CLK(dco_clk),
    .D(_01947_),
    .Q( execution_unit_0.register_file_0.r4_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09184_ (
    .CLK(dco_clk),
    .D(_01948_),
    .Q( execution_unit_0.register_file_0.r4_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09185_ (
    .CLK(dco_clk),
    .D(_01949_),
    .Q( execution_unit_0.register_file_0.r4_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09186_ (
    .CLK(dco_clk),
    .D(_01950_),
    .Q( execution_unit_0.register_file_0.r4_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09187_ (
    .CLK(dco_clk),
    .D(_01951_),
    .Q( execution_unit_0.register_file_0.r4_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09188_ (
    .CLK(dco_clk),
    .D(_01952_),
    .Q( execution_unit_0.register_file_0.r4_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09189_ (
    .CLK(dco_clk),
    .D(_01953_),
    .Q( execution_unit_0.register_file_0.r4_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09190_ (
    .CLK(dco_clk),
    .D(_01954_),
    .Q( execution_unit_0.register_file_0.r4_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09191_ (
    .CLK(dco_clk),
    .D(_01955_),
    .Q( execution_unit_0.register_file_0.r3_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09192_ (
    .CLK(dco_clk),
    .D(_01956_),
    .Q( execution_unit_0.register_file_0.r3_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09193_ (
    .CLK(dco_clk),
    .D(_01957_),
    .Q( execution_unit_0.register_file_0.r3_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09194_ (
    .CLK(dco_clk),
    .D(_01958_),
    .Q( execution_unit_0.register_file_0.r3_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09195_ (
    .CLK(dco_clk),
    .D(_01959_),
    .Q( execution_unit_0.register_file_0.r3_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09196_ (
    .CLK(dco_clk),
    .D(_01960_),
    .Q( execution_unit_0.register_file_0.r3_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09197_ (
    .CLK(dco_clk),
    .D(_01961_),
    .Q( execution_unit_0.register_file_0.r3_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09198_ (
    .CLK(dco_clk),
    .D(_01962_),
    .Q( execution_unit_0.register_file_0.r3_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09199_ (
    .CLK(dco_clk),
    .D(_01963_),
    .Q( execution_unit_0.register_file_0.r3_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09200_ (
    .CLK(dco_clk),
    .D(_01964_),
    .Q( execution_unit_0.register_file_0.r3_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09201_ (
    .CLK(dco_clk),
    .D(_01965_),
    .Q( execution_unit_0.register_file_0.r3_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09202_ (
    .CLK(dco_clk),
    .D(_01966_),
    .Q( execution_unit_0.register_file_0.r3_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09203_ (
    .CLK(dco_clk),
    .D(_01967_),
    .Q( execution_unit_0.register_file_0.r3_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09204_ (
    .CLK(dco_clk),
    .D(_01968_),
    .Q( execution_unit_0.register_file_0.r3_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09205_ (
    .CLK(dco_clk),
    .D(_01969_),
    .Q( execution_unit_0.register_file_0.r3_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09206_ (
    .CLK(dco_clk),
    .D(_01970_),
    .Q( execution_unit_0.register_file_0.r3_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09207_ (
    .CLK(dco_clk),
    .D(_01971_),
    .Q( execution_unit_0.alu_0.status_0_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09208_ (
    .CLK(dco_clk),
    .D(_01755_),
    .Q( execution_unit_0.register_file_0.r2_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09209_ (
    .CLK(dco_clk),
    .D(_01972_),
    .Q( execution_unit_0.register_file_0.r1_1_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09210_ (
    .CLK(dco_clk),
    .D(_01973_),
    .Q( execution_unit_0.register_file_0.r1_2_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09211_ (
    .CLK(dco_clk),
    .D(_01974_),
    .Q( execution_unit_0.register_file_0.r1_3_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09212_ (
    .CLK(dco_clk),
    .D(_01975_),
    .Q( execution_unit_0.register_file_0.r1_4_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09213_ (
    .CLK(dco_clk),
    .D(_01976_),
    .Q( execution_unit_0.register_file_0.r1_5_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09214_ (
    .CLK(dco_clk),
    .D(_01977_),
    .Q( execution_unit_0.register_file_0.r1_6_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09215_ (
    .CLK(dco_clk),
    .D(_01978_),
    .Q( execution_unit_0.register_file_0.r1_7_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09216_ (
    .CLK(dco_clk),
    .D(_01979_),
    .Q( execution_unit_0.register_file_0.r1_8_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09217_ (
    .CLK(dco_clk),
    .D(_01980_),
    .Q( execution_unit_0.register_file_0.r1_9_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09218_ (
    .CLK(dco_clk),
    .D(_01981_),
    .Q( execution_unit_0.register_file_0.r1_10_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09219_ (
    .CLK(dco_clk),
    .D(_01982_),
    .Q( execution_unit_0.register_file_0.r1_11_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09220_ (
    .CLK(dco_clk),
    .D(_01983_),
    .Q( execution_unit_0.register_file_0.r1_12_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09221_ (
    .CLK(dco_clk),
    .D(_01984_),
    .Q( execution_unit_0.register_file_0.r1_13_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09222_ (
    .CLK(dco_clk),
    .D(_01985_),
    .Q( execution_unit_0.register_file_0.r1_14_ ),
    .R(_01756_),
    .S(1'h1)
  );
  DFFSR _09223_ (
    .CLK(dco_clk),
    .D(_01986_),
    .Q( execution_unit_0.register_file_0.r1_15_ ),
    .R(_01756_),
    .S(1'h1)
  );
  INVX1 _09224_ (
    .A(cpu_en),
    .Y(_03167_)
  );
  INVX1 _09225_ (
    .A( frontend_0.i_state_1_ ),
    .Y(_03168_)
  );
  INVX1 _09226_ (
    .A( frontend_0.i_state_0_ ),
    .Y(_03169_)
  );
  INVX1 _09227_ (
    .A( frontend_0.i_state_2_ ),
    .Y(_03170_)
  );
  INVX1 _09228_ (
    .A(irq_5_),
    .Y(_03171_)
  );
  INVX1 _09229_ (
    .A(irq_7_),
    .Y(_03172_)
  );
  INVX1 _09230_ (
    .A(irq_9_),
    .Y(_03173_)
  );
  INVX1 _09231_ (
    .A(irq_11_),
    .Y(_03174_)
  );
  INVX1 _09232_ (
    .A(irq_12_),
    .Y(_03175_)
  );
  INVX1 _09233_ (
    .A( execution_unit_0.gie ),
    .Y(_03176_)
  );
  INVX1 _09234_ (
    .A(1'h0),
    .Y(_03177_)
  );
  INVX1 _09235_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_03178_)
  );
  INVX1 _09236_ (
    .A( frontend_0.exec_jmp ),
    .Y(_03179_)
  );
  INVX1 _09237_ (
    .A( frontend_0.exec_dst_wr ),
    .Y(_03180_)
  );
  INVX1 _09238_ (
    .A( frontend_0.exec_src_wr ),
    .Y(_03181_)
  );
  INVX1 _09239_ (
    .A( execution_unit_0.e_state_1_ ),
    .Y(_03182_)
  );
  INVX1 _09240_ (
    .A( execution_unit_0.e_state_2_ ),
    .Y(_03183_)
  );
  INVX1 _09241_ (
    .A( execution_unit_0.e_state_3_ ),
    .Y(_03184_)
  );
  INVX1 _09242_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .Y(_03185_)
  );
  INVX1 _09243_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .Y(_03186_)
  );
  INVX1 _09244_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .Y(_03187_)
  );
  INVX1 _09245_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .Y(_03188_)
  );
  INVX1 _09246_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .Y(_03189_)
  );
  INVX1 _09247_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .Y(_03190_)
  );
  INVX1 _09248_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .Y(_03191_)
  );
  INVX1 _09249_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .Y(_03192_)
  );
  INVX1 _09250_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .Y(_03193_)
  );
  INVX1 _09251_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .Y(_03194_)
  );
  INVX1 _09252_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .Y(_03195_)
  );
  INVX1 _09253_ (
    .A( execution_unit_0.inst_as_4_ ),
    .Y(_03196_)
  );
  INVX1 _09254_ (
    .A( frontend_0.exec_dext_rdy ),
    .Y(_03197_)
  );
  INVX1 _09255_ (
    .A( execution_unit_0.UNUSED_inst_ad_idx ),
    .Y(_03198_)
  );
  INVX1 _09256_ (
    .A( execution_unit_0.pc_sw_wr ),
    .Y(_03199_)
  );
  INVX1 _09257_ (
    .A( frontend_0.inst_sz_1_ ),
    .Y(_03200_)
  );
  INVX1 _09258_ (
    .A( execution_unit_0.inst_type_0_ ),
    .Y(_03201_)
  );
  INVX1 _09259_ (
    .A( execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_03202_)
  );
  INVX1 _09260_ (
    .A( dbg_0.UNUSED_pc_1_ ),
    .Y(_03203_)
  );
  INVX1 _09261_ (
    .A( frontend_0.irq_addr_1_ ),
    .Y(_03204_)
  );
  INVX1 _09262_ (
    .A( dbg_0.UNUSED_pc_2_ ),
    .Y(_03205_)
  );
  INVX1 _09263_ (
    .A( frontend_0.irq_addr_2_ ),
    .Y(_03206_)
  );
  INVX1 _09264_ (
    .A( dbg_0.UNUSED_pc_3_ ),
    .Y(_03207_)
  );
  INVX1 _09265_ (
    .A( frontend_0.irq_addr_3_ ),
    .Y(_03208_)
  );
  INVX1 _09266_ (
    .A( dbg_0.UNUSED_pc_4_ ),
    .Y(_03209_)
  );
  INVX1 _09267_ (
    .A( dbg_0.UNUSED_pc_5_ ),
    .Y(_03210_)
  );
  INVX1 _09268_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .Y(_03211_)
  );
  INVX1 _09269_ (
    .A( dbg_0.UNUSED_pc_7_ ),
    .Y(_03212_)
  );
  INVX1 _09270_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .Y(_03213_)
  );
  INVX1 _09271_ (
    .A( dbg_0.UNUSED_pc_9_ ),
    .Y(_03214_)
  );
  INVX1 _09272_ (
    .A( dbg_0.UNUSED_pc_10_ ),
    .Y(_03215_)
  );
  INVX1 _09273_ (
    .A( dbg_0.UNUSED_pc_11_ ),
    .Y(_03216_)
  );
  INVX1 _09274_ (
    .A( dbg_0.UNUSED_pc_12_ ),
    .Y(_03217_)
  );
  INVX1 _09275_ (
    .A( dbg_0.UNUSED_pc_13_ ),
    .Y(_03218_)
  );
  INVX1 _09276_ (
    .A( dbg_0.UNUSED_pc_14_ ),
    .Y(_03219_)
  );
  INVX1 _09277_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .Y(_03220_)
  );
  INVX1 _09278_ (
    .A( frontend_0.inst_dest_bin_2_ ),
    .Y(_03221_)
  );
  INVX1 _09279_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .Y(_03222_)
  );
  INVX1 _09280_ (
    .A( execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_03223_)
  );
  INVX1 _09281_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .Y(_03224_)
  );
  INVX1 _09282_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .Y(_03225_)
  );
  INVX1 _09283_ (
    .A( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03226_)
  );
  INVX1 _09284_ (
    .A( frontend_0.inst_jmp_bin_1_ ),
    .Y(_03227_)
  );
  INVX1 _09285_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .Y(_03228_)
  );
  INVX1 _09286_ (
    .A( frontend_0.inst_src_bin_1_ ),
    .Y(_03229_)
  );
  INVX1 _09287_ (
    .A( frontend_0.inst_src_bin_0_ ),
    .Y(_03230_)
  );
  INVX1 _09288_ (
    .A( execution_unit_0.inst_type_2_ ),
    .Y(_03231_)
  );
  INVX1 _09289_ (
    .A( frontend_0.pmem_busy ),
    .Y(_03232_)
  );
  INVX1 _09290_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .Y(_03233_)
  );
  INVX1 _09291_ (
    .A(_05695_),
    .Y(_02907_)
  );
  INVX1 _09292_ (
    .A( execution_unit_0.inst_dext_14_ ),
    .Y(_03234_)
  );
  INVX1 _09293_ (
    .A( execution_unit_0.inst_sext_2_ ),
    .Y(_03235_)
  );
  INVX1 _09294_ (
    .A( execution_unit_0.inst_sext_4_ ),
    .Y(_03236_)
  );
  INVX1 _09295_ (
    .A( execution_unit_0.inst_sext_5_ ),
    .Y(_03237_)
  );
  INVX1 _09296_ (
    .A( execution_unit_0.inst_sext_6_ ),
    .Y(_03238_)
  );
  INVX1 _09297_ (
    .A( execution_unit_0.inst_sext_7_ ),
    .Y(_03239_)
  );
  INVX1 _09298_ (
    .A( execution_unit_0.inst_sext_8_ ),
    .Y(_03240_)
  );
  INVX1 _09299_ (
    .A( execution_unit_0.inst_sext_9_ ),
    .Y(_03241_)
  );
  INVX1 _09300_ (
    .A( execution_unit_0.inst_sext_10_ ),
    .Y(_03242_)
  );
  INVX1 _09301_ (
    .A( execution_unit_0.inst_sext_11_ ),
    .Y(_03243_)
  );
  INVX1 _09302_ (
    .A( execution_unit_0.inst_sext_12_ ),
    .Y(_03244_)
  );
  INVX1 _09303_ (
    .A( execution_unit_0.inst_sext_13_ ),
    .Y(_03245_)
  );
  INVX1 _09304_ (
    .A( execution_unit_0.inst_sext_14_ ),
    .Y(_03246_)
  );
  INVX1 _09305_ (
    .A( execution_unit_0.inst_sext_15_ ),
    .Y(_03247_)
  );
  INVX1 _09306_ (
    .A( execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_03248_)
  );
  INVX1 _09307_ (
    .A( execution_unit_0.inst_as_7_ ),
    .Y(_03249_)
  );
  NOR2X1 _09308_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03250_)
  );
  OR2X1 _09309_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03251_)
  );
  NAND2X1 _09310_ (
    .A( execution_unit_0.e_state_2_ ),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_03252_)
  );
  OAI21X1 _09311_ (
    .A(_03251_),
    .B(_03252_),
    .C( frontend_0.exec_jmp ),
    .Y(_03253_)
  );
  NAND2X1 _09312_ (
    .A(_03183_),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_03254_)
  );
  OR2X1 _09313_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03182_),
    .Y(_03255_)
  );
  NOR2X1 _09314_ (
    .A(_03254_),
    .B(_03255_),
    .Y(_03256_)
  );
  OR2X1 _09315_ (
    .A(_03254_),
    .B(_03255_),
    .Y(_03257_)
  );
  OAI21X1 _09316_ (
    .A(_03254_),
    .B(_03255_),
    .C( frontend_0.exec_dst_wr ),
    .Y(_03258_)
  );
  AND2X1 _09317_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03259_)
  );
  NAND2X1 _09318_ (
    .A( execution_unit_0.e_state_0_ ),
    .B( execution_unit_0.e_state_1_ ),
    .Y(_03260_)
  );
  NAND2X1 _09319_ (
    .A( execution_unit_0.e_state_2_ ),
    .B(_03184_),
    .Y(_03261_)
  );
  NOR3X1 _09320_ (
    .A(_03183_),
    .B( execution_unit_0.e_state_3_ ),
    .C(_03260_),
    .Y(_03262_)
  );
  NAND3X1 _09321_ (
    .A(_03183_),
    .B( execution_unit_0.e_state_3_ ),
    .C(_03259_),
    .Y(_03263_)
  );
  NOR2X1 _09322_ (
    .A( frontend_0.exec_src_wr ),
    .B(_03263_),
    .Y(_03264_)
  );
  OR2X1 _09323_ (
    .A( frontend_0.exec_src_wr ),
    .B(_03263_),
    .Y(_03265_)
  );
  AOI21X1 _09324_ (
    .A( frontend_0.exec_src_wr ),
    .B(_03262_),
    .C( frontend_0.exec_dst_wr ),
    .Y(_03266_)
  );
  AOI22X1 _09325_ (
    .A( frontend_0.exec_dst_wr ),
    .B(_03257_),
    .C(_03265_),
    .D(_03266_),
    .Y(_03267_)
  );
  OAI21X1 _09326_ (
    .A( frontend_0.exec_jmp ),
    .B(_03267_),
    .C(_03253_),
    .Y(_03268_)
  );
  INVX1 _09327_ (
    .A(_03268_),
    .Y( execution_unit_0.exec_done )
  );
  NOR2X1 _09328_ (
    .A( frontend_0.i_state_1_ ),
    .B(_03169_),
    .Y(_03269_)
  );
  NAND2X1 _09329_ (
    .A(_03168_),
    .B( frontend_0.i_state_0_ ),
    .Y(_03270_)
  );
  NOR2X1 _09330_ (
    .A(_03170_),
    .B(_03270_),
    .Y(_03271_)
  );
  NAND2X1 _09331_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03269_),
    .Y(_03272_)
  );
  NOR3X1 _09332_ (
    .A(irq_11_),
    .B(irq_10_),
    .C( frontend_0.wdt_irq ),
    .Y(_03273_)
  );
  NOR2X1 _09333_ (
    .A(irq_9_),
    .B(irq_8_),
    .Y(_03274_)
  );
  NAND2X1 _09334_ (
    .A(_03273_),
    .B(_03274_),
    .Y(_03275_)
  );
  NOR2X1 _09335_ (
    .A(irq_5_),
    .B(irq_4_),
    .Y(_03276_)
  );
  NOR2X1 _09336_ (
    .A(irq_3_),
    .B(irq_2_),
    .Y(_03277_)
  );
  NAND2X1 _09337_ (
    .A(_03276_),
    .B(_03277_),
    .Y(_03278_)
  );
  NOR2X1 _09338_ (
    .A(irq_7_),
    .B(irq_6_),
    .Y(_03279_)
  );
  NOR2X1 _09339_ (
    .A(irq_13_),
    .B(irq_12_),
    .Y(_03280_)
  );
  OR2X1 _09340_ (
    .A(irq_13_),
    .B(irq_12_),
    .Y(_03281_)
  );
  NOR2X1 _09341_ (
    .A(irq_1_),
    .B(irq_0_),
    .Y(_03282_)
  );
  NAND3X1 _09342_ (
    .A(_03279_),
    .B(_03280_),
    .C(_03282_),
    .Y(_03283_)
  );
  NOR3X1 _09343_ (
    .A(_03275_),
    .B(_03278_),
    .C(_03283_),
    .Y(_03284_)
  );
  OAI21X1 _09344_ (
    .A(_03176_),
    .B(_03284_),
    .C(_03177_),
    .Y(_03285_)
  );
  OR2X1 _09345_ (
    .A( dbg_0.dbg_halt_cmd ),
    .B(_03167_),
    .Y(_03286_)
  );
  NOR2X1 _09346_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_03286_),
    .Y(_03287_)
  );
  AND2X1 _09347_ (
    .A(_03285_),
    .B(_03287_),
    .Y(_03288_)
  );
  NAND2X1 _09348_ (
    .A(_03285_),
    .B(_03287_),
    .Y(_03289_)
  );
  AOI21X1 _09349_ (
    .A(_03268_),
    .B(_03272_),
    .C(_03289_),
    .Y(_03290_)
  );
  OAI21X1 _09350_ (
    .A( execution_unit_0.exec_done ),
    .B(_03271_),
    .C(_03288_),
    .Y(_03291_)
  );
  NOR2X1 _09351_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.fe_mdb_in_15_ ),
    .Y(_03292_)
  );
  INVX1 _09352_ (
    .A(_03292_),
    .Y(_03293_)
  );
  NOR3X1 _09353_ (
    .A(_03186_),
    .B(_03290_),
    .C(_03293_),
    .Y(_03294_)
  );
  NAND3X1 _09354_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03291_),
    .C(_03292_),
    .Y(_03295_)
  );
  NAND2X1 _09355_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03295_),
    .Y(_03296_)
  );
  NAND3X1 _09356_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B( dbg_0.fe_mdb_in_4_ ),
    .C(_03295_),
    .Y(_03297_)
  );
  INVX1 _09357_ (
    .A(_03297_),
    .Y(_03298_)
  );
  NAND3X1 _09358_ (
    .A(_03186_),
    .B(_03291_),
    .C(_03292_),
    .Y(_03299_)
  );
  INVX1 _09359_ (
    .A(_03299_),
    .Y(_03300_)
  );
  NOR2X1 _09360_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B( dbg_0.fe_mdb_in_3_ ),
    .Y(_03301_)
  );
  NAND2X1 _09361_ (
    .A(_03188_),
    .B(_03189_),
    .Y(_03302_)
  );
  NOR2X1 _09362_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B( dbg_0.fe_mdb_in_11_ ),
    .Y(_03303_)
  );
  INVX1 _09363_ (
    .A(_03303_),
    .Y(_03304_)
  );
  MUX2X1 _09364_ (
    .A(_03304_),
    .B(_03302_),
    .S(_03299_),
    .Y(_03305_)
  );
  MUX2X1 _09365_ (
    .A(_03303_),
    .B(_03301_),
    .S(_03299_),
    .Y(_03306_)
  );
  MUX2X1 _09366_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B( dbg_0.fe_mdb_in_0_ ),
    .S(_03299_),
    .Y(_03307_)
  );
  MUX2X1 _09367_ (
    .A(_03190_),
    .B(_03191_),
    .S(_03299_),
    .Y(_03308_)
  );
  MUX2X1 _09368_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B( dbg_0.fe_mdb_in_1_ ),
    .S(_03299_),
    .Y(_03309_)
  );
  MUX2X1 _09369_ (
    .A(_03192_),
    .B(_03193_),
    .S(_03299_),
    .Y(_03310_)
  );
  NAND2X1 _09370_ (
    .A(_03305_),
    .B(_03310_),
    .Y(_03311_)
  );
  AOI21X1 _09371_ (
    .A(_03308_),
    .B(_03309_),
    .C(_03306_),
    .Y(_03312_)
  );
  NOR2X1 _09372_ (
    .A(_03297_),
    .B(_03312_),
    .Y(_03313_)
  );
  OR2X1 _09373_ (
    .A(_03297_),
    .B(_03312_),
    .Y(_03314_)
  );
  NOR3X1 _09374_ (
    .A(_03306_),
    .B(_03308_),
    .C(_03310_),
    .Y(_03315_)
  );
  NAND3X1 _09375_ (
    .A(_03305_),
    .B(_03307_),
    .C(_03309_),
    .Y(_03316_)
  );
  NOR2X1 _09376_ (
    .A(_03297_),
    .B(_03316_),
    .Y(_03317_)
  );
  NAND2X1 _09377_ (
    .A(_03298_),
    .B(_03315_),
    .Y(_03318_)
  );
  NAND2X1 _09378_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03195_),
    .Y(_03319_)
  );
  NOR2X1 _09379_ (
    .A(_03192_),
    .B(_03299_),
    .Y(_03320_)
  );
  OR2X1 _09380_ (
    .A(_03192_),
    .B(_03299_),
    .Y(_03321_)
  );
  OR2X1 _09381_ (
    .A(_03319_),
    .B(_03321_),
    .Y(_03322_)
  );
  NOR3X1 _09382_ (
    .A(_03194_),
    .B( dbg_0.fe_mdb_in_4_ ),
    .C(_03294_),
    .Y(_03323_)
  );
  OAI21X1 _09383_ (
    .A(_03306_),
    .B(_03309_),
    .C(_03323_),
    .Y(_03324_)
  );
  AND2X1 _09384_ (
    .A(_03322_),
    .B(_03324_),
    .Y(_03325_)
  );
  OAI21X1 _09385_ (
    .A(_03319_),
    .B(_03321_),
    .C(_03324_),
    .Y(_03326_)
  );
  NOR3X1 _09386_ (
    .A(_03313_),
    .B(_03317_),
    .C(_03326_),
    .Y(_03327_)
  );
  NAND3X1 _09387_ (
    .A(_03314_),
    .B(_03318_),
    .C(_03325_),
    .Y(_03328_)
  );
  NOR2X1 _09388_ (
    .A(_03290_),
    .B(_03292_),
    .Y(_03329_)
  );
  AND2X1 _09389_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03329_),
    .Y(_03330_)
  );
  NAND2X1 _09390_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03329_),
    .Y(_03331_)
  );
  NOR2X1 _09391_ (
    .A( clock_module_0.UNUSED_cpuoff ),
    .B(_03286_),
    .Y(_03332_)
  );
  OR2X1 _09392_ (
    .A( clock_module_0.UNUSED_cpuoff ),
    .B(_03286_),
    .Y(_03333_)
  );
  NOR2X1 _09393_ (
    .A(_03271_),
    .B(_03333_),
    .Y(_03334_)
  );
  OAI21X1 _09394_ (
    .A(_03170_),
    .B(_03270_),
    .C(_03332_),
    .Y(_03335_)
  );
  NOR3X1 _09395_ (
    .A(_03306_),
    .B(_03307_),
    .C(_03309_),
    .Y(_03336_)
  );
  NAND3X1 _09396_ (
    .A(_03305_),
    .B(_03308_),
    .C(_03310_),
    .Y(_03337_)
  );
  NAND2X1 _09397_ (
    .A(_03194_),
    .B( dbg_0.fe_mdb_in_4_ ),
    .Y(_03338_)
  );
  NOR2X1 _09398_ (
    .A(_03294_),
    .B(_03338_),
    .Y(_03339_)
  );
  OR2X1 _09399_ (
    .A(_03294_),
    .B(_03338_),
    .Y(_03340_)
  );
  AOI21X1 _09400_ (
    .A(_03337_),
    .B(_03339_),
    .C(_03335_),
    .Y(_03341_)
  );
  OAI21X1 _09401_ (
    .A(_03336_),
    .B(_03340_),
    .C(_03334_),
    .Y(_03342_)
  );
  OAI21X1 _09402_ (
    .A(_03328_),
    .B(_03330_),
    .C(_03341_),
    .Y(_03343_)
  );
  NOR2X1 _09403_ (
    .A( frontend_0.exec_dst_wr ),
    .B(_03263_),
    .Y(_03344_)
  );
  AND2X1 _09404_ (
    .A(_03179_),
    .B(_03344_),
    .Y(_03345_)
  );
  INVX1 _09405_ (
    .A(_03345_),
    .Y(_03346_)
  );
  NOR2X1 _09406_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_03252_),
    .Y(_03347_)
  );
  NOR2X1 _09407_ (
    .A(_03262_),
    .B(_03347_),
    .Y(_03348_)
  );
  OAI21X1 _09408_ (
    .A(_03254_),
    .B(_03255_),
    .C(_03348_),
    .Y(_03349_)
  );
  NAND2X1 _09409_ (
    .A( frontend_0.exec_jmp ),
    .B(_03348_),
    .Y(_03350_)
  );
  NAND2X1 _09410_ (
    .A(_03349_),
    .B(_03350_),
    .Y(_03351_)
  );
  NAND2X1 _09411_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B( dbg_0.fe_mdb_in_7_ ),
    .Y(_03352_)
  );
  OR2X1 _09412_ (
    .A(_03321_),
    .B(_03352_),
    .Y(_03353_)
  );
  OAI21X1 _09413_ (
    .A(_03321_),
    .B(_03352_),
    .C(_03291_),
    .Y(_03354_)
  );
  NAND2X1 _09414_ (
    .A(_03178_),
    .B(_03354_),
    .Y(_03355_)
  );
  AND2X1 _09415_ (
    .A(_03178_),
    .B(_03354_),
    .Y(_03356_)
  );
  AOI21X1 _09416_ (
    .A(_03346_),
    .B(_03351_),
    .C(_03356_),
    .Y(_03357_)
  );
  NOR2X1 _09417_ (
    .A(_03251_),
    .B(_03254_),
    .Y(_03358_)
  );
  NOR2X1 _09418_ (
    .A(_03168_),
    .B( frontend_0.i_state_2_ ),
    .Y(_03359_)
  );
  NAND2X1 _09419_ (
    .A( frontend_0.i_state_0_ ),
    .B(_03359_),
    .Y(_03360_)
  );
  INVX1 _09420_ (
    .A(_03360_),
    .Y(_03361_)
  );
  NOR2X1 _09421_ (
    .A( execution_unit_0.inst_as_1_ ),
    .B( execution_unit_0.inst_as_4_ ),
    .Y(_03362_)
  );
  NOR2X1 _09422_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B( execution_unit_0.inst_as_5_ ),
    .Y(_03363_)
  );
  NAND2X1 _09423_ (
    .A(_03362_),
    .B(_03363_),
    .Y(_03364_)
  );
  NOR2X1 _09424_ (
    .A(_03360_),
    .B(_03364_),
    .Y(_03365_)
  );
  NOR2X1 _09425_ (
    .A( frontend_0.i_state_1_ ),
    .B( frontend_0.i_state_0_ ),
    .Y(_03366_)
  );
  NAND2X1 _09426_ (
    .A(_03168_),
    .B(_03169_),
    .Y(_03367_)
  );
  AOI21X1 _09427_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03366_),
    .C(_03365_),
    .Y(_03368_)
  );
  INVX1 _09428_ (
    .A(_03368_),
    .Y(_03369_)
  );
  OAI21X1 _09429_ (
    .A( frontend_0.exec_dext_rdy ),
    .B(_03369_),
    .C(_03358_),
    .Y(_03370_)
  );
  NAND2X1 _09430_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03182_),
    .Y(_03371_)
  );
  OR2X1 _09431_ (
    .A(_03261_),
    .B(_03371_),
    .Y(_03372_)
  );
  INVX1 _09432_ (
    .A(_03372_),
    .Y(_03373_)
  );
  NAND2X1 _09433_ (
    .A(_03361_),
    .B(_03364_),
    .Y(_03374_)
  );
  NOR2X1 _09434_ (
    .A(_03255_),
    .B(_03261_),
    .Y(_03375_)
  );
  NOR2X1 _09435_ (
    .A( execution_unit_0.UNUSED_inst_ad_symb ),
    .B( execution_unit_0.inst_ad_6_ ),
    .Y(_03376_)
  );
  NAND3X1 _09436_ (
    .A(_03198_),
    .B(_03375_),
    .C(_03376_),
    .Y(_03377_)
  );
  NOR2X1 _09437_ (
    .A(_03254_),
    .B(_03371_),
    .Y(_03378_)
  );
  INVX1 _09438_ (
    .A(_03378_),
    .Y(_03379_)
  );
  OAI21X1 _09439_ (
    .A(_03251_),
    .B(_03261_),
    .C(_03379_),
    .Y(_03380_)
  );
  NOR2X1 _09440_ (
    .A( execution_unit_0.e_state_2_ ),
    .B( execution_unit_0.e_state_3_ ),
    .Y(_03381_)
  );
  INVX1 _09441_ (
    .A(_03381_),
    .Y(_03382_)
  );
  OAI21X1 _09442_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03382_),
    .C(_03377_),
    .Y(_03383_)
  );
  NOR2X1 _09443_ (
    .A(_03380_),
    .B(_03383_),
    .Y(_03384_)
  );
  AOI22X1 _09444_ (
    .A( frontend_0.exec_src_wr ),
    .B(_03345_),
    .C(_03373_),
    .D(_03374_),
    .Y(_03385_)
  );
  NAND3X1 _09445_ (
    .A(_03370_),
    .B(_03384_),
    .C(_03385_),
    .Y(_03386_)
  );
  AOI21X1 _09446_ (
    .A(_03343_),
    .B(_03357_),
    .C(_03386_),
    .Y(_03387_)
  );
  INVX1 _09447_ (
    .A(_03387_),
    .Y( frontend_0.e_state_nxt_0_ )
  );
  AOI22X1 _09448_ (
    .A(_03298_),
    .B(_03315_),
    .C(_03337_),
    .D(_03339_),
    .Y(_03388_)
  );
  OAI22X1 _09449_ (
    .A(_03297_),
    .B(_03316_),
    .C(_03336_),
    .D(_03340_),
    .Y(_03389_)
  );
  NOR3X1 _09450_ (
    .A(_03313_),
    .B(_03326_),
    .C(_03389_),
    .Y(_03390_)
  );
  NAND3X1 _09451_ (
    .A(_03314_),
    .B(_03325_),
    .C(_03388_),
    .Y(_03391_)
  );
  NOR2X1 _09452_ (
    .A(_03344_),
    .B(_03349_),
    .Y(_03392_)
  );
  NOR2X1 _09453_ (
    .A(_03356_),
    .B(_03392_),
    .Y(_03393_)
  );
  OAI21X1 _09454_ (
    .A(_03344_),
    .B(_03349_),
    .C(_03355_),
    .Y(_03394_)
  );
  AOI21X1 _09455_ (
    .A(_03327_),
    .B(_03341_),
    .C(_03394_),
    .Y(_03395_)
  );
  OAI21X1 _09456_ (
    .A(_03328_),
    .B(_03342_),
    .C(_03393_),
    .Y(_03396_)
  );
  NAND2X1 _09457_ (
    .A( frontend_0.exec_jmp ),
    .B(_03256_),
    .Y(_03397_)
  );
  AOI21X1 _09458_ (
    .A(_03259_),
    .B(_03381_),
    .C(_03373_),
    .Y(_03398_)
  );
  OAI21X1 _09459_ (
    .A(_03179_),
    .B(_03257_),
    .C(_03398_),
    .Y(_03399_)
  );
  INVX1 _09460_ (
    .A(_03399_),
    .Y(_03400_)
  );
  OAI21X1 _09461_ (
    .A( frontend_0.exec_jmp ),
    .B( frontend_0.exec_src_wr ),
    .C(_03344_),
    .Y(_03401_)
  );
  AND2X1 _09462_ (
    .A(_03400_),
    .B(_03401_),
    .Y(_03402_)
  );
  NAND2X1 _09463_ (
    .A(_03400_),
    .B(_03401_),
    .Y(_03403_)
  );
  NAND2X1 _09464_ (
    .A(_03396_),
    .B(_03402_),
    .Y( frontend_0.e_state_nxt_2_ )
  );
  NOR2X1 _09465_ (
    .A(_03264_),
    .B(_03349_),
    .Y(_03404_)
  );
  NOR2X1 _09466_ (
    .A(_03356_),
    .B(_03404_),
    .Y(_03405_)
  );
  OAI21X1 _09467_ (
    .A(_03264_),
    .B(_03349_),
    .C(_03355_),
    .Y(_03406_)
  );
  AOI21X1 _09468_ (
    .A(_03334_),
    .B(_03391_),
    .C(_03406_),
    .Y(_03407_)
  );
  OAI21X1 _09469_ (
    .A(_03335_),
    .B(_03390_),
    .C(_03405_),
    .Y(_03408_)
  );
  AOI22X1 _09470_ (
    .A(_03179_),
    .B(_03180_),
    .C(_03263_),
    .D(_03397_),
    .Y(_03409_)
  );
  OAI22X1 _09471_ (
    .A( execution_unit_0.e_state_1_ ),
    .B(_03254_),
    .C(_03261_),
    .D( execution_unit_0.e_state_0_ ),
    .Y(_03410_)
  );
  NOR2X1 _09472_ (
    .A(_03409_),
    .B(_03410_),
    .Y(_03411_)
  );
  INVX1 _09473_ (
    .A(_03411_),
    .Y(_03412_)
  );
  NAND2X1 _09474_ (
    .A(_03408_),
    .B(_03411_),
    .Y( frontend_0.e_state_nxt_3_ )
  );
  NAND2X1 _09475_ (
    .A(_03331_),
    .B(_03388_),
    .Y(_03413_)
  );
  INVX1 _09476_ (
    .A(_03413_),
    .Y(_03414_)
  );
  AND2X1 _09477_ (
    .A(_03169_),
    .B(_03359_),
    .Y(_03415_)
  );
  OAI21X1 _09478_ (
    .A(_03252_),
    .B(_03371_),
    .C(_03268_),
    .Y(_03416_)
  );
  INVX1 _09479_ (
    .A(_03416_),
    .Y(_03417_)
  );
  NAND2X1 _09480_ (
    .A(_03415_),
    .B(_03416_),
    .Y(_03418_)
  );
  INVX1 _09481_ (
    .A(_03418_),
    .Y( dbg_0.decode_noirq )
  );
  AND2X1 _09482_ (
    .A(_03291_),
    .B(_03415_),
    .Y(_03419_)
  );
  NOR2X1 _09483_ (
    .A(_03290_),
    .B(_03418_),
    .Y(_03420_)
  );
  NAND2X1 _09484_ (
    .A(_03291_),
    .B( dbg_0.decode_noirq ),
    .Y(_03421_)
  );
  NAND3X1 _09485_ (
    .A(_03199_),
    .B(_03413_),
    .C(_03420_),
    .Y(_03422_)
  );
  NOR2X1 _09486_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03367_),
    .Y(_03423_)
  );
  NAND2X1 _09487_ (
    .A(_03170_),
    .B(_03366_),
    .Y(_03424_)
  );
  NOR2X1 _09488_ (
    .A(_03272_),
    .B(_03332_),
    .Y(_03425_)
  );
  NAND3X1 _09489_ (
    .A( execution_unit_0.e_state_0_ ),
    .B(_03286_),
    .C(_03347_),
    .Y(_03426_)
  );
  AOI21X1 _09490_ (
    .A(_03268_),
    .B(_03426_),
    .C(_03332_),
    .Y(_03427_)
  );
  AOI22X1 _09491_ (
    .A(_03289_),
    .B(_03425_),
    .C(_03427_),
    .D(_03419_),
    .Y(_03428_)
  );
  AND2X1 _09492_ (
    .A(_03424_),
    .B(_03428_),
    .Y(_03429_)
  );
  NAND2X1 _09493_ (
    .A(_03422_),
    .B(_03429_),
    .Y( frontend_0.i_state_nxt_0_ )
  );
  AOI21X1 _09494_ (
    .A( frontend_0.inst_sz_0_ ),
    .B(_03200_),
    .C( execution_unit_0.pc_sw_wr ),
    .Y(_03430_)
  );
  INVX1 _09495_ (
    .A(_03430_),
    .Y(_03431_)
  );
  OAI21X1 _09496_ (
    .A(_03360_),
    .B(_03431_),
    .C(_03428_),
    .Y( frontend_0.i_state_nxt_2_ )
  );
  NOR2X1 _09497_ (
    .A(_03272_),
    .B(_03333_),
    .Y(_03432_)
  );
  OAI21X1 _09498_ (
    .A(_03415_),
    .B(_03432_),
    .C(_03291_),
    .Y(_03433_)
  );
  NAND2X1 _09499_ (
    .A(_03361_),
    .B(_03431_),
    .Y(_03434_)
  );
  NOR2X1 _09500_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03270_),
    .Y(_03435_)
  );
  NAND2X1 _09501_ (
    .A(_03170_),
    .B(_03269_),
    .Y(_03436_)
  );
  OAI21X1 _09502_ (
    .A(_03360_),
    .B(_03430_),
    .C(_03436_),
    .Y(_03437_)
  );
  AOI21X1 _09503_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03366_),
    .C(_03437_),
    .Y(_03438_)
  );
  OAI21X1 _09504_ (
    .A(_03427_),
    .B(_03433_),
    .C(_03438_),
    .Y( frontend_0.i_state_nxt_1_ )
  );
  OAI21X1 _09505_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03321_),
    .C(_03331_),
    .Y(_03439_)
  );
  AOI21X1 _09506_ (
    .A(_03327_),
    .B(_03439_),
    .C(_03342_),
    .Y(_03440_)
  );
  NOR2X1 _09507_ (
    .A(_03356_),
    .B(_03440_),
    .Y(_03441_)
  );
  AOI21X1 _09508_ (
    .A(_03181_),
    .B(_03441_),
    .C( frontend_0.exec_jmp ),
    .Y(_03442_)
  );
  NOR2X1 _09509_ (
    .A( frontend_0.exec_dst_wr ),
    .B(_03442_),
    .Y(_03443_)
  );
  NOR2X1 _09510_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .Y(_03444_)
  );
  NOR2X1 _09511_ (
    .A(_03182_),
    .B(_03252_),
    .Y(_03445_)
  );
  NOR2X1 _09512_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_03377_),
    .Y(_03446_)
  );
  AOI21X1 _09513_ (
    .A(_03184_),
    .B(_03250_),
    .C(_03378_),
    .Y(_03447_)
  );
  OAI21X1 _09514_ (
    .A(_03372_),
    .B(_03374_),
    .C(_03447_),
    .Y(_03448_)
  );
  AOI21X1 _09515_ (
    .A(_03444_),
    .B(_03446_),
    .C(_03448_),
    .Y(_03449_)
  );
  OAI21X1 _09516_ (
    .A(_03351_),
    .B(_03441_),
    .C(_03449_),
    .Y(_03450_)
  );
  NOR2X1 _09517_ (
    .A(_03445_),
    .B(_03450_),
    .Y(_03451_)
  );
  OAI21X1 _09518_ (
    .A(_03263_),
    .B(_03443_),
    .C(_03451_),
    .Y( frontend_0.e_state_nxt_1_ )
  );
  OAI21X1 _09519_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03367_),
    .C(_03199_),
    .Y(_03452_)
  );
  AOI21X1 _09520_ (
    .A(_03191_),
    .B(_03435_),
    .C(_03452_),
    .Y(_03453_)
  );
  OAI21X1 _09521_ (
    .A( dbg_0.UNUSED_pc_0_ ),
    .B(_03435_),
    .C(_03453_),
    .Y(_03454_)
  );
  OAI21X1 _09522_ (
    .A(_03199_),
    .B(_03202_),
    .C(_03454_),
    .Y( execution_unit_0.pc_nxt_0_ )
  );
  NOR2X1 _09523_ (
    .A(_03199_),
    .B( execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_03455_)
  );
  NAND2X1 _09524_ (
    .A(_03415_),
    .B(_03417_),
    .Y(_03456_)
  );
  AOI22X1 _09525_ (
    .A(_03396_),
    .B(_03402_),
    .C(_03408_),
    .D(_03411_),
    .Y(_03457_)
  );
  OAI22X1 _09526_ (
    .A(_03395_),
    .B(_03403_),
    .C(_03407_),
    .D(_03412_),
    .Y(_03458_)
  );
  AOI22X1 _09527_ (
    .A(_03415_),
    .B(_03417_),
    .C(_03457_),
    .D( frontend_0.e_state_nxt_0_ ),
    .Y(_03459_)
  );
  OAI21X1 _09528_ (
    .A(_03387_),
    .B(_03458_),
    .C(_03456_),
    .Y(_03460_)
  );
  XNOR2X1 _09529_ (
    .A(_03203_),
    .B(_03459_),
    .Y(_03461_)
  );
  AOI21X1 _09530_ (
    .A(_03193_),
    .B(_03435_),
    .C(_03423_),
    .Y(_03462_)
  );
  OAI21X1 _09531_ (
    .A(_03435_),
    .B(_03461_),
    .C(_03462_),
    .Y(_03463_)
  );
  AOI21X1 _09532_ (
    .A( frontend_0.irq_addr_1_ ),
    .B(_03423_),
    .C( execution_unit_0.pc_sw_wr ),
    .Y(_03464_)
  );
  AOI21X1 _09533_ (
    .A(_03463_),
    .B(_03464_),
    .C(_03455_),
    .Y( execution_unit_0.pc_nxt_1_ )
  );
  NOR2X1 _09534_ (
    .A(_03199_),
    .B( execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_03465_)
  );
  OAI21X1 _09535_ (
    .A(_03203_),
    .B(_03460_),
    .C(_03205_),
    .Y(_03466_)
  );
  NOR3X1 _09536_ (
    .A(_03203_),
    .B(_03205_),
    .C(_03460_),
    .Y(_03467_)
  );
  NAND3X1 _09537_ (
    .A( dbg_0.UNUSED_pc_1_ ),
    .B( dbg_0.UNUSED_pc_2_ ),
    .C(_03459_),
    .Y(_03468_)
  );
  AOI21X1 _09538_ (
    .A(_03466_),
    .B(_03468_),
    .C(_03435_),
    .Y(_03469_)
  );
  OAI21X1 _09539_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B(_03436_),
    .C(_03424_),
    .Y(_03470_)
  );
  OR2X1 _09540_ (
    .A(_03469_),
    .B(_03470_),
    .Y(_03471_)
  );
  AOI21X1 _09541_ (
    .A( frontend_0.irq_addr_2_ ),
    .B(_03423_),
    .C( execution_unit_0.pc_sw_wr ),
    .Y(_03472_)
  );
  AOI21X1 _09542_ (
    .A(_03471_),
    .B(_03472_),
    .C(_03465_),
    .Y( execution_unit_0.pc_nxt_2_ )
  );
  NOR2X1 _09543_ (
    .A(_03199_),
    .B( execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_03473_)
  );
  XNOR2X1 _09544_ (
    .A(_03207_),
    .B(_03467_),
    .Y(_03474_)
  );
  NOR2X1 _09545_ (
    .A(_03435_),
    .B(_03474_),
    .Y(_03475_)
  );
  OAI21X1 _09546_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .B(_03436_),
    .C(_03424_),
    .Y(_03476_)
  );
  NAND2X1 _09547_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03423_),
    .Y(_03477_)
  );
  OAI21X1 _09548_ (
    .A(_03475_),
    .B(_03476_),
    .C(_03477_),
    .Y(_03478_)
  );
  NOR2X1 _09549_ (
    .A( execution_unit_0.pc_sw_wr ),
    .B(_03478_),
    .Y(_03479_)
  );
  NOR2X1 _09550_ (
    .A(_03473_),
    .B(_03479_),
    .Y( execution_unit_0.pc_nxt_3_ )
  );
  OAI21X1 _09551_ (
    .A(_03207_),
    .B(_03468_),
    .C(_03209_),
    .Y(_03480_)
  );
  NOR3X1 _09552_ (
    .A(_03207_),
    .B(_03209_),
    .C(_03468_),
    .Y(_03481_)
  );
  NAND3X1 _09553_ (
    .A( dbg_0.UNUSED_pc_3_ ),
    .B( dbg_0.UNUSED_pc_4_ ),
    .C(_03467_),
    .Y(_03482_)
  );
  AOI21X1 _09554_ (
    .A(_03480_),
    .B(_03482_),
    .C(_03435_),
    .Y(_03483_)
  );
  OAI21X1 _09555_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03436_),
    .C(_03424_),
    .Y(_03484_)
  );
  NAND2X1 _09556_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03423_),
    .Y(_03485_)
  );
  OAI21X1 _09557_ (
    .A(_03483_),
    .B(_03484_),
    .C(_03485_),
    .Y(_03486_)
  );
  MUX2X1 _09558_ (
    .A( execution_unit_0.alu_0.alu_out_4_ ),
    .B(_03486_),
    .S( execution_unit_0.pc_sw_wr ),
    .Y(_03487_)
  );
  INVX1 _09559_ (
    .A(_03487_),
    .Y( execution_unit_0.pc_nxt_4_ )
  );
  NOR2X1 _09560_ (
    .A(_03210_),
    .B(_03482_),
    .Y(_03488_)
  );
  OAI21X1 _09561_ (
    .A( dbg_0.UNUSED_pc_5_ ),
    .B(_03481_),
    .C(_03436_),
    .Y(_03489_)
  );
  AOI21X1 _09562_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03490_)
  );
  OAI21X1 _09563_ (
    .A(_03488_),
    .B(_03489_),
    .C(_03490_),
    .Y(_03491_)
  );
  OAI21X1 _09564_ (
    .A(_03199_),
    .B( execution_unit_0.alu_0.alu_out_5_ ),
    .C(_03491_),
    .Y(_03492_)
  );
  INVX1 _09565_ (
    .A(_03492_),
    .Y( execution_unit_0.pc_nxt_5_ )
  );
  NOR3X1 _09566_ (
    .A(_03210_),
    .B(_03211_),
    .C(_03482_),
    .Y(_03493_)
  );
  NAND3X1 _09567_ (
    .A( dbg_0.UNUSED_pc_5_ ),
    .B( dbg_0.UNUSED_pc_6_ ),
    .C(_03481_),
    .Y(_03494_)
  );
  OAI21X1 _09568_ (
    .A( dbg_0.UNUSED_pc_6_ ),
    .B(_03488_),
    .C(_03436_),
    .Y(_03495_)
  );
  AOI21X1 _09569_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03496_)
  );
  OAI21X1 _09570_ (
    .A(_03493_),
    .B(_03495_),
    .C(_03496_),
    .Y(_03497_)
  );
  OAI21X1 _09571_ (
    .A(_03199_),
    .B( execution_unit_0.alu_0.alu_out_6_ ),
    .C(_03497_),
    .Y(_03498_)
  );
  INVX1 _09572_ (
    .A(_03498_),
    .Y( execution_unit_0.pc_nxt_6_ )
  );
  NOR2X1 _09573_ (
    .A(_03212_),
    .B(_03494_),
    .Y(_03499_)
  );
  OAI21X1 _09574_ (
    .A( dbg_0.UNUSED_pc_7_ ),
    .B(_03493_),
    .C(_03436_),
    .Y(_03500_)
  );
  AOI21X1 _09575_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03501_)
  );
  OAI21X1 _09576_ (
    .A(_03499_),
    .B(_03500_),
    .C(_03501_),
    .Y(_03502_)
  );
  OAI21X1 _09577_ (
    .A(_03199_),
    .B( execution_unit_0.alu_0.alu_out_7_ ),
    .C(_03502_),
    .Y(_03503_)
  );
  INVX1 _09578_ (
    .A(_03503_),
    .Y( execution_unit_0.pc_nxt_7_ )
  );
  NOR3X1 _09579_ (
    .A(_03212_),
    .B(_03213_),
    .C(_03494_),
    .Y(_03504_)
  );
  NAND3X1 _09580_ (
    .A( dbg_0.UNUSED_pc_7_ ),
    .B( dbg_0.UNUSED_pc_8_ ),
    .C(_03493_),
    .Y(_03505_)
  );
  OAI21X1 _09581_ (
    .A( dbg_0.UNUSED_pc_8_ ),
    .B(_03499_),
    .C(_03436_),
    .Y(_03506_)
  );
  AOI21X1 _09582_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03507_)
  );
  OAI21X1 _09583_ (
    .A(_03504_),
    .B(_03506_),
    .C(_03507_),
    .Y(_03508_)
  );
  OAI21X1 _09584_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_8_ ),
    .C(_03508_),
    .Y(_03509_)
  );
  INVX1 _09585_ (
    .A(_03509_),
    .Y( execution_unit_0.pc_nxt_8_ )
  );
  NOR2X1 _09586_ (
    .A(_03214_),
    .B(_03505_),
    .Y(_03510_)
  );
  OAI21X1 _09587_ (
    .A( dbg_0.UNUSED_pc_9_ ),
    .B(_03504_),
    .C(_03436_),
    .Y(_03511_)
  );
  AOI21X1 _09588_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03512_)
  );
  OAI21X1 _09589_ (
    .A(_03510_),
    .B(_03511_),
    .C(_03512_),
    .Y(_03513_)
  );
  OAI21X1 _09590_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_9_ ),
    .C(_03513_),
    .Y(_03514_)
  );
  INVX1 _09591_ (
    .A(_03514_),
    .Y( execution_unit_0.pc_nxt_9_ )
  );
  NOR3X1 _09592_ (
    .A(_03214_),
    .B(_03215_),
    .C(_03505_),
    .Y(_03515_)
  );
  NAND3X1 _09593_ (
    .A( dbg_0.UNUSED_pc_9_ ),
    .B( dbg_0.UNUSED_pc_10_ ),
    .C(_03504_),
    .Y(_03516_)
  );
  OAI21X1 _09594_ (
    .A( dbg_0.UNUSED_pc_10_ ),
    .B(_03510_),
    .C(_03436_),
    .Y(_03517_)
  );
  AOI21X1 _09595_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03518_)
  );
  OAI21X1 _09596_ (
    .A(_03515_),
    .B(_03517_),
    .C(_03518_),
    .Y(_03519_)
  );
  OAI21X1 _09597_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_10_ ),
    .C(_03519_),
    .Y(_03520_)
  );
  INVX1 _09598_ (
    .A(_03520_),
    .Y( execution_unit_0.pc_nxt_10_ )
  );
  XNOR2X1 _09599_ (
    .A( dbg_0.UNUSED_pc_11_ ),
    .B(_03515_),
    .Y(_03521_)
  );
  AOI21X1 _09600_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03522_)
  );
  OAI21X1 _09601_ (
    .A(_03435_),
    .B(_03521_),
    .C(_03522_),
    .Y(_03523_)
  );
  OAI21X1 _09602_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_11_ ),
    .C(_03523_),
    .Y(_03524_)
  );
  INVX1 _09603_ (
    .A(_03524_),
    .Y( execution_unit_0.pc_nxt_11_ )
  );
  NAND3X1 _09604_ (
    .A( dbg_0.UNUSED_pc_11_ ),
    .B( dbg_0.UNUSED_pc_12_ ),
    .C(_03515_),
    .Y(_03525_)
  );
  OAI21X1 _09605_ (
    .A(_03216_),
    .B(_03516_),
    .C(_03217_),
    .Y(_03526_)
  );
  NAND2X1 _09606_ (
    .A(_03525_),
    .B(_03526_),
    .Y(_03527_)
  );
  AOI21X1 _09607_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03528_)
  );
  OAI21X1 _09608_ (
    .A(_03435_),
    .B(_03527_),
    .C(_03528_),
    .Y(_03529_)
  );
  OAI21X1 _09609_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_12_ ),
    .C(_03529_),
    .Y(_03530_)
  );
  INVX1 _09610_ (
    .A(_03530_),
    .Y( execution_unit_0.pc_nxt_12_ )
  );
  XNOR2X1 _09611_ (
    .A(_03218_),
    .B(_03525_),
    .Y(_03531_)
  );
  AOI21X1 _09612_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03532_)
  );
  OAI21X1 _09613_ (
    .A(_03435_),
    .B(_03531_),
    .C(_03532_),
    .Y(_03533_)
  );
  OAI21X1 _09614_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_13_ ),
    .C(_03533_),
    .Y(_03534_)
  );
  INVX1 _09615_ (
    .A(_03534_),
    .Y( execution_unit_0.pc_nxt_13_ )
  );
  NOR2X1 _09616_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_14_ ),
    .Y(_03535_)
  );
  NOR3X1 _09617_ (
    .A(_03218_),
    .B(_03219_),
    .C(_03525_),
    .Y(_03536_)
  );
  OAI21X1 _09618_ (
    .A(_03218_),
    .B(_03525_),
    .C(_03219_),
    .Y(_03537_)
  );
  OAI21X1 _09619_ (
    .A( frontend_0.i_state_2_ ),
    .B(_03270_),
    .C(_03537_),
    .Y(_03538_)
  );
  OR2X1 _09620_ (
    .A(_03536_),
    .B(_03538_),
    .Y(_03539_)
  );
  AOI21X1 _09621_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03540_)
  );
  AOI21X1 _09622_ (
    .A(_03539_),
    .B(_03540_),
    .C(_03535_),
    .Y( execution_unit_0.pc_nxt_14_ )
  );
  OR2X1 _09623_ (
    .A(_03199_),
    .B( execution_unit_0.pc_sw_15_ ),
    .Y(_03541_)
  );
  XNOR2X1 _09624_ (
    .A( dbg_0.UNUSED_pc_15_ ),
    .B(_03536_),
    .Y(_03542_)
  );
  AOI21X1 _09625_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03435_),
    .C(_03452_),
    .Y(_03543_)
  );
  OAI21X1 _09626_ (
    .A(_03435_),
    .B(_03542_),
    .C(_03543_),
    .Y(_03544_)
  );
  AND2X1 _09627_ (
    .A(_03541_),
    .B(_03544_),
    .Y( execution_unit_0.pc_nxt_15_ )
  );
  NOR2X1 _09628_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03545_)
  );
  NAND2X1 _09629_ (
    .A(_03221_),
    .B(_03545_),
    .Y(_03546_)
  );
  OR2X1 _09630_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03546_),
    .Y(_03547_)
  );
  NAND2X1 _09631_ (
    .A(_03223_),
    .B(_03444_),
    .Y(_03548_)
  );
  NOR2X1 _09632_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B( execution_unit_0.inst_type_1_ ),
    .Y(_03549_)
  );
  OAI21X1 _09633_ (
    .A(_03547_),
    .B(_03548_),
    .C(_03549_),
    .Y(_03550_)
  );
  NAND2X1 _09634_ (
    .A(_03225_),
    .B(_03226_),
    .Y(_03551_)
  );
  OR2X1 _09635_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_03551_),
    .Y(_03552_)
  );
  OAI21X1 _09636_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_03552_),
    .C( dbg_0.cpu_stat_full_0_ ),
    .Y(_03553_)
  );
  AND2X1 _09637_ (
    .A(_03550_),
    .B(_03553_),
    .Y( execution_unit_0.inst_dest_0_ )
  );
  AND2X1 _09638_ (
    .A(_03222_),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03554_)
  );
  NAND2X1 _09639_ (
    .A(_03221_),
    .B(_03554_),
    .Y(_03555_)
  );
  NOR2X1 _09640_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03555_),
    .Y(_03556_)
  );
  OAI21X1 _09641_ (
    .A(_03548_),
    .B(_03556_),
    .C(_03549_),
    .Y(_03557_)
  );
  NAND3X1 _09642_ (
    .A(_03224_),
    .B(_03225_),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03558_)
  );
  XOR2X1 _09643_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .B(_03552_),
    .Y(_03559_)
  );
  NAND2X1 _09644_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .B(_03559_),
    .Y(_03560_)
  );
  OAI21X1 _09645_ (
    .A(_03558_),
    .B(_03560_),
    .C(_03557_),
    .Y( execution_unit_0.inst_dest_1_ )
  );
  NOR2X1 _09646_ (
    .A(_03222_),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03561_)
  );
  NAND2X1 _09647_ (
    .A(_03221_),
    .B(_03561_),
    .Y(_03562_)
  );
  OR2X1 _09648_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03562_),
    .Y(_03563_)
  );
  NAND3X1 _09649_ (
    .A(_03223_),
    .B(_03444_),
    .C(_03549_),
    .Y(_03564_)
  );
  NAND3X1 _09650_ (
    .A(_03224_),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C(_03226_),
    .Y(_03565_)
  );
  OAI22X1 _09651_ (
    .A(_03563_),
    .B(_03564_),
    .C(_03565_),
    .D(_03560_),
    .Y( execution_unit_0.inst_dest_2_ )
  );
  NAND2X1 _09652_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .B( frontend_0.inst_dest_bin_0_ ),
    .Y(_03566_)
  );
  NOR2X1 _09653_ (
    .A( frontend_0.inst_dest_bin_2_ ),
    .B(_03566_),
    .Y(_03567_)
  );
  NAND2X1 _09654_ (
    .A(_03220_),
    .B(_03567_),
    .Y(_03568_)
  );
  NAND3X1 _09655_ (
    .A(_03224_),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03569_)
  );
  OAI22X1 _09656_ (
    .A(_03564_),
    .B(_03568_),
    .C(_03569_),
    .D(_03560_),
    .Y( execution_unit_0.inst_dest_3_ )
  );
  NAND3X1 _09657_ (
    .A(_03220_),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03545_),
    .Y(_03570_)
  );
  OR2X1 _09658_ (
    .A(_03224_),
    .B(_03551_),
    .Y(_03571_)
  );
  OAI22X1 _09659_ (
    .A(_03564_),
    .B(_03570_),
    .C(_03571_),
    .D(_03560_),
    .Y( execution_unit_0.inst_dest_4_ )
  );
  NAND3X1 _09660_ (
    .A(_03220_),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03554_),
    .Y(_03572_)
  );
  NAND3X1 _09661_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B(_03225_),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03573_)
  );
  OAI22X1 _09662_ (
    .A(_03564_),
    .B(_03572_),
    .C(_03573_),
    .D(_03560_),
    .Y( execution_unit_0.inst_dest_5_ )
  );
  NAND3X1 _09663_ (
    .A(_03220_),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03561_),
    .Y(_03574_)
  );
  NAND3X1 _09664_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C(_03226_),
    .Y(_03575_)
  );
  OAI22X1 _09665_ (
    .A(_03564_),
    .B(_03574_),
    .C(_03575_),
    .D(_03560_),
    .Y( execution_unit_0.inst_dest_6_ )
  );
  OR2X1 _09666_ (
    .A(_03221_),
    .B(_03566_),
    .Y(_03576_)
  );
  OR2X1 _09667_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03576_),
    .Y(_03577_)
  );
  NAND3X1 _09668_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .B( dbg_0.dbg_mem_addr_1_ ),
    .C( dbg_0.dbg_mem_addr_0_ ),
    .Y(_03578_)
  );
  OAI22X1 _09669_ (
    .A(_03564_),
    .B(_03577_),
    .C(_03578_),
    .D(_03560_),
    .Y( execution_unit_0.inst_dest_7_ )
  );
  OR2X1 _09670_ (
    .A(_03220_),
    .B(_03546_),
    .Y(_03579_)
  );
  OAI22X1 _09671_ (
    .A(_03552_),
    .B(_03553_),
    .C(_03564_),
    .D(_03579_),
    .Y( execution_unit_0.inst_dest_8_ )
  );
  OR2X1 _09672_ (
    .A(_03220_),
    .B(_03555_),
    .Y(_03580_)
  );
  OR2X1 _09673_ (
    .A(_03178_),
    .B(_03559_),
    .Y(_03581_)
  );
  OAI22X1 _09674_ (
    .A(_03564_),
    .B(_03580_),
    .C(_03581_),
    .D(_03558_),
    .Y( execution_unit_0.inst_dest_9_ )
  );
  OR2X1 _09675_ (
    .A(_03220_),
    .B(_03562_),
    .Y(_03582_)
  );
  OAI22X1 _09676_ (
    .A(_03565_),
    .B(_03581_),
    .C(_03582_),
    .D(_03564_),
    .Y( execution_unit_0.inst_dest_10_ )
  );
  NAND2X1 _09677_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03567_),
    .Y(_03583_)
  );
  OAI22X1 _09678_ (
    .A(_03569_),
    .B(_03581_),
    .C(_03583_),
    .D(_03564_),
    .Y( execution_unit_0.inst_dest_11_ )
  );
  NAND3X1 _09679_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03545_),
    .Y(_03584_)
  );
  OAI22X1 _09680_ (
    .A(_03571_),
    .B(_03581_),
    .C(_03584_),
    .D(_03564_),
    .Y( execution_unit_0.inst_dest_12_ )
  );
  NAND3X1 _09681_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03554_),
    .Y(_03585_)
  );
  OAI22X1 _09682_ (
    .A(_03573_),
    .B(_03581_),
    .C(_03585_),
    .D(_03564_),
    .Y( execution_unit_0.inst_dest_13_ )
  );
  NAND3X1 _09683_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B( frontend_0.inst_dest_bin_2_ ),
    .C(_03561_),
    .Y(_03586_)
  );
  OAI22X1 _09684_ (
    .A(_03575_),
    .B(_03581_),
    .C(_03586_),
    .D(_03564_),
    .Y( execution_unit_0.inst_dest_14_ )
  );
  OR2X1 _09685_ (
    .A(_03220_),
    .B(_03576_),
    .Y(_03587_)
  );
  OAI22X1 _09686_ (
    .A(_03578_),
    .B(_03581_),
    .C(_03587_),
    .D(_03564_),
    .Y( execution_unit_0.inst_dest_15_ )
  );
  OAI21X1 _09687_ (
    .A(_03201_),
    .B(_03547_),
    .C(_03223_),
    .Y(_03588_)
  );
  NOR2X1 _09688_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B( execution_unit_0.inst_type_2_ ),
    .Y(_03589_)
  );
  NAND2X1 _09689_ (
    .A(_03588_),
    .B(_03589_),
    .Y(_03590_)
  );
  NAND2X1 _09690_ (
    .A(_03229_),
    .B(_03230_),
    .Y(_03591_)
  );
  OR2X1 _09691_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B(_03591_),
    .Y(_03592_)
  );
  OR2X1 _09692_ (
    .A( frontend_0.inst_jmp_bin_1_ ),
    .B(_03592_),
    .Y(_03593_)
  );
  OAI21X1 _09693_ (
    .A(_03231_),
    .B(_03593_),
    .C(_03590_),
    .Y( execution_unit_0.inst_src_0_ )
  );
  NOR2X1 _09694_ (
    .A(_03201_),
    .B( execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_03594_)
  );
  AOI21X1 _09695_ (
    .A(_03556_),
    .B(_03594_),
    .C( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_03595_)
  );
  NAND3X1 _09696_ (
    .A(_03228_),
    .B(_03229_),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03596_)
  );
  XNOR2X1 _09697_ (
    .A(_03227_),
    .B(_03592_),
    .Y(_03597_)
  );
  NAND2X1 _09698_ (
    .A( execution_unit_0.inst_type_2_ ),
    .B(_03597_),
    .Y(_03598_)
  );
  OAI22X1 _09699_ (
    .A( execution_unit_0.inst_type_2_ ),
    .B(_03595_),
    .C(_03596_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_1_ )
  );
  NAND2X1 _09700_ (
    .A(_03589_),
    .B(_03594_),
    .Y(_03599_)
  );
  NAND3X1 _09701_ (
    .A(_03228_),
    .B( frontend_0.inst_src_bin_1_ ),
    .C(_03230_),
    .Y(_03600_)
  );
  OAI22X1 _09702_ (
    .A(_03563_),
    .B(_03599_),
    .C(_03600_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_2_ )
  );
  NAND3X1 _09703_ (
    .A(_03228_),
    .B( frontend_0.inst_src_bin_1_ ),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03601_)
  );
  OAI22X1 _09704_ (
    .A(_03568_),
    .B(_03599_),
    .C(_03601_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_3_ )
  );
  OR2X1 _09705_ (
    .A(_03228_),
    .B(_03591_),
    .Y(_03602_)
  );
  OAI22X1 _09706_ (
    .A(_03570_),
    .B(_03599_),
    .C(_03602_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_4_ )
  );
  NAND3X1 _09707_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B(_03229_),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03603_)
  );
  OAI22X1 _09708_ (
    .A(_03572_),
    .B(_03599_),
    .C(_03603_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_5_ )
  );
  NAND3X1 _09709_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B( frontend_0.inst_src_bin_1_ ),
    .C(_03230_),
    .Y(_03604_)
  );
  OAI22X1 _09710_ (
    .A(_03574_),
    .B(_03599_),
    .C(_03604_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_6_ )
  );
  NAND3X1 _09711_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B( frontend_0.inst_src_bin_1_ ),
    .C( frontend_0.inst_src_bin_0_ ),
    .Y(_03605_)
  );
  OAI22X1 _09712_ (
    .A(_03577_),
    .B(_03599_),
    .C(_03605_),
    .D(_03598_),
    .Y( execution_unit_0.inst_src_7_ )
  );
  NAND2X1 _09713_ (
    .A( frontend_0.inst_jmp_bin_1_ ),
    .B( execution_unit_0.inst_type_2_ ),
    .Y(_03606_)
  );
  OAI22X1 _09714_ (
    .A(_03579_),
    .B(_03599_),
    .C(_03606_),
    .D(_03592_),
    .Y( execution_unit_0.inst_src_8_ )
  );
  OR2X1 _09715_ (
    .A(_03231_),
    .B(_03597_),
    .Y(_03607_)
  );
  OAI22X1 _09716_ (
    .A(_03580_),
    .B(_03599_),
    .C(_03607_),
    .D(_03596_),
    .Y( execution_unit_0.inst_src_9_ )
  );
  OAI22X1 _09717_ (
    .A(_03582_),
    .B(_03599_),
    .C(_03600_),
    .D(_03607_),
    .Y( execution_unit_0.inst_src_10_ )
  );
  OAI22X1 _09718_ (
    .A(_03583_),
    .B(_03599_),
    .C(_03601_),
    .D(_03607_),
    .Y( execution_unit_0.inst_src_11_ )
  );
  OAI22X1 _09719_ (
    .A(_03584_),
    .B(_03599_),
    .C(_03602_),
    .D(_03607_),
    .Y( execution_unit_0.inst_src_12_ )
  );
  OAI22X1 _09720_ (
    .A(_03585_),
    .B(_03599_),
    .C(_03603_),
    .D(_03607_),
    .Y( execution_unit_0.inst_src_13_ )
  );
  OAI22X1 _09721_ (
    .A(_03586_),
    .B(_03599_),
    .C(_03604_),
    .D(_03607_),
    .Y( execution_unit_0.inst_src_14_ )
  );
  OAI22X1 _09722_ (
    .A(_03587_),
    .B(_03599_),
    .C(_03605_),
    .D(_03607_),
    .Y( execution_unit_0.inst_src_15_ )
  );
  NAND2X1 _09723_ (
    .A(_03204_),
    .B(_03206_),
    .Y(_03608_)
  );
  OR2X1 _09724_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03608_),
    .Y(_03609_)
  );
  OR2X1 _09725_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03609_),
    .Y(_03610_)
  );
  NOR2X1 _09726_ (
    .A(_03424_),
    .B(_03610_),
    .Y(_05616_)
  );
  NAND3X1 _09727_ (
    .A( frontend_0.irq_addr_1_ ),
    .B(_03206_),
    .C(_03208_),
    .Y(_03611_)
  );
  XOR2X1 _09728_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03609_),
    .Y(_03612_)
  );
  NAND2X1 _09729_ (
    .A(_03423_),
    .B(_03612_),
    .Y(_03613_)
  );
  NOR2X1 _09730_ (
    .A(_03611_),
    .B(_03613_),
    .Y(_05621_)
  );
  NAND3X1 _09731_ (
    .A(_03204_),
    .B( frontend_0.irq_addr_2_ ),
    .C(_03208_),
    .Y(_03614_)
  );
  NOR2X1 _09732_ (
    .A(_03613_),
    .B(_03614_),
    .Y(_05622_)
  );
  NAND2X1 _09733_ (
    .A( frontend_0.irq_addr_1_ ),
    .B( frontend_0.irq_addr_2_ ),
    .Y(_03615_)
  );
  OR2X1 _09734_ (
    .A( frontend_0.irq_addr_3_ ),
    .B(_03615_),
    .Y(_03616_)
  );
  NOR2X1 _09735_ (
    .A(_03613_),
    .B(_03616_),
    .Y(_05623_)
  );
  OR2X1 _09736_ (
    .A(_03208_),
    .B(_03608_),
    .Y(_03617_)
  );
  NOR2X1 _09737_ (
    .A(_03613_),
    .B(_03617_),
    .Y(_05624_)
  );
  NAND3X1 _09738_ (
    .A( frontend_0.irq_addr_1_ ),
    .B(_03206_),
    .C( frontend_0.irq_addr_3_ ),
    .Y(_03618_)
  );
  NOR2X1 _09739_ (
    .A(_03613_),
    .B(_03618_),
    .Y(_05625_)
  );
  NAND3X1 _09740_ (
    .A(_03204_),
    .B( frontend_0.irq_addr_2_ ),
    .C( frontend_0.irq_addr_3_ ),
    .Y(_03619_)
  );
  NOR2X1 _09741_ (
    .A(_03613_),
    .B(_03619_),
    .Y(_05626_)
  );
  NOR2X1 _09742_ (
    .A(_03477_),
    .B(_03615_),
    .Y(_03620_)
  );
  AND2X1 _09743_ (
    .A(_03612_),
    .B(_03620_),
    .Y(_05627_)
  );
  NOR2X1 _09744_ (
    .A(_03485_),
    .B(_03609_),
    .Y(_05628_)
  );
  OR2X1 _09745_ (
    .A(_03424_),
    .B(_03612_),
    .Y(_03621_)
  );
  NOR2X1 _09746_ (
    .A(_03611_),
    .B(_03621_),
    .Y(_05629_)
  );
  NOR2X1 _09747_ (
    .A(_03614_),
    .B(_03621_),
    .Y(_05617_)
  );
  NOR2X1 _09748_ (
    .A(_03616_),
    .B(_03621_),
    .Y(_05618_)
  );
  NOR2X1 _09749_ (
    .A(_03485_),
    .B(_03617_),
    .Y(_05619_)
  );
  NOR2X1 _09750_ (
    .A(_03618_),
    .B(_03621_),
    .Y(_05620_)
  );
  OAI21X1 _09751_ (
    .A(_03178_),
    .B(_03286_),
    .C(_03232_),
    .Y(_03622_)
  );
  NOR2X1 _09752_ (
    .A(_03452_),
    .B(_03622_),
    .Y(_03623_)
  );
  NAND2X1 _09753_ (
    .A(_03460_),
    .B(_03623_),
    .Y( frontend_0.mb_en )
  );
  NAND2X1 _09754_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_03227_),
    .Y(_03624_)
  );
  OR2X1 _09755_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B(_03624_),
    .Y(_03625_)
  );
  NOR2X1 _09756_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B(_03625_),
    .Y( execution_unit_0.alu_0.inst_jmp_0_ )
  );
  OR2X1 _09757_ (
    .A(_03228_),
    .B(_03624_),
    .Y(_03626_)
  );
  NOR2X1 _09758_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B(_03626_),
    .Y( execution_unit_0.alu_0.inst_jmp_1_ )
  );
  NAND2X1 _09759_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .Y(_03627_)
  );
  OR2X1 _09760_ (
    .A( frontend_0.inst_jmp_bin_0_ ),
    .B(_03627_),
    .Y(_03628_)
  );
  NOR2X1 _09761_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B(_03628_),
    .Y( execution_unit_0.alu_0.inst_jmp_2_ )
  );
  OR2X1 _09762_ (
    .A(_03228_),
    .B(_03627_),
    .Y(_03629_)
  );
  NOR2X1 _09763_ (
    .A( frontend_0.inst_jmp_bin_2_ ),
    .B(_03629_),
    .Y( execution_unit_0.alu_0.inst_jmp_3_ )
  );
  NOR2X1 _09764_ (
    .A(_03233_),
    .B(_03625_),
    .Y( execution_unit_0.alu_0.inst_jmp_4_ )
  );
  NOR2X1 _09765_ (
    .A(_03233_),
    .B(_03626_),
    .Y( execution_unit_0.alu_0.inst_jmp_5_ )
  );
  NOR2X1 _09766_ (
    .A(_03233_),
    .B(_03628_),
    .Y( execution_unit_0.alu_0.inst_jmp_6_ )
  );
  OAI21X1 _09767_ (
    .A( dbg_0.dbg_halt_cmd ),
    .B(_03167_),
    .C( frontend_0.i_state_nxt_2_ ),
    .Y(_03630_)
  );
  AOI21X1 _09768_ (
    .A(_03422_),
    .B(_03429_),
    .C(_03630_),
    .Y(_02906_)
  );
  AOI21X1 _09769_ (
    .A(_03197_),
    .B(_03368_),
    .C(_03378_),
    .Y(_02920_)
  );
  NAND2X1 _09770_ (
    .A( execution_unit_0.inst_type_0_ ),
    .B(_03375_),
    .Y(_03631_)
  );
  OAI21X1 _09771_ (
    .A(_03260_),
    .B(_03261_),
    .C( frontend_0.exec_src_wr ),
    .Y(_03632_)
  );
  OAI21X1 _09772_ (
    .A(_03256_),
    .B(_03632_),
    .C(_03631_),
    .Y(_02921_)
  );
  OAI21X1 _09773_ (
    .A(_03254_),
    .B(_03371_),
    .C(_03258_),
    .Y(_02922_)
  );
  AND2X1 _09774_ (
    .A(_03295_),
    .B(_03322_),
    .Y(_03633_)
  );
  NOR2X1 _09775_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_03302_),
    .Y(_03634_)
  );
  NAND3X1 _09776_ (
    .A(_03193_),
    .B(_03329_),
    .C(_03634_),
    .Y(_03635_)
  );
  OAI21X1 _09777_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03635_),
    .C(_03633_),
    .Y(_03636_)
  );
  INVX1 _09778_ (
    .A(_03636_),
    .Y(_03637_)
  );
  NOR2X1 _09779_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .Y(_03638_)
  );
  NAND2X1 _09780_ (
    .A(_03291_),
    .B(_03418_),
    .Y(_03639_)
  );
  OAI21X1 _09781_ (
    .A(_03637_),
    .B(_03638_),
    .C(_03253_),
    .Y(_02923_)
  );
  MUX2X1 _09782_ (
    .A( execution_unit_0.inst_dext_0_ ),
    .B( dbg_0.fe_mdb_in_0_ ),
    .S(_03368_),
    .Y(_03640_)
  );
  INVX1 _09783_ (
    .A(_03640_),
    .Y(_02955_)
  );
  OAI22X1 _09784_ (
    .A(_03170_),
    .B(_03367_),
    .C(_03434_),
    .D( execution_unit_0.inst_as_4_ ),
    .Y(_03641_)
  );
  NAND2X1 _09785_ (
    .A( execution_unit_0.UNUSED_inst_ad_symb ),
    .B(_03641_),
    .Y(_03642_)
  );
  OAI21X1 _09786_ (
    .A(_03196_),
    .B(_03360_),
    .C(_03642_),
    .Y(_03643_)
  );
  AND2X1 _09787_ (
    .A(_03193_),
    .B(_03643_),
    .Y(_03644_)
  );
  NOR2X1 _09788_ (
    .A(_03193_),
    .B(_03643_),
    .Y(_03645_)
  );
  NOR2X1 _09789_ (
    .A(_03644_),
    .B(_03645_),
    .Y(_03646_)
  );
  NAND2X1 _09790_ (
    .A( execution_unit_0.inst_dext_1_ ),
    .B(_03368_),
    .Y(_03647_)
  );
  OAI21X1 _09791_ (
    .A(_03368_),
    .B(_03646_),
    .C(_03647_),
    .Y(_02956_)
  );
  XNOR2X1 _09792_ (
    .A( dbg_0.fe_mdb_in_2_ ),
    .B(_03644_),
    .Y(_03648_)
  );
  NAND2X1 _09793_ (
    .A( execution_unit_0.inst_dext_2_ ),
    .B(_03368_),
    .Y(_03649_)
  );
  OAI21X1 _09794_ (
    .A(_03368_),
    .B(_03648_),
    .C(_03649_),
    .Y(_02957_)
  );
  AOI21X1 _09795_ (
    .A(_03188_),
    .B(_03644_),
    .C(_03189_),
    .Y(_03650_)
  );
  NAND2X1 _09796_ (
    .A(_03301_),
    .B(_03644_),
    .Y(_03651_)
  );
  AOI21X1 _09797_ (
    .A(_03301_),
    .B(_03644_),
    .C(_03650_),
    .Y(_03652_)
  );
  NAND2X1 _09798_ (
    .A( execution_unit_0.inst_dext_3_ ),
    .B(_03368_),
    .Y(_03653_)
  );
  OAI21X1 _09799_ (
    .A(_03368_),
    .B(_03652_),
    .C(_03653_),
    .Y(_02958_)
  );
  XOR2X1 _09800_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03651_),
    .Y(_03654_)
  );
  NAND2X1 _09801_ (
    .A( execution_unit_0.inst_dext_4_ ),
    .B(_03368_),
    .Y(_03655_)
  );
  OAI21X1 _09802_ (
    .A(_03368_),
    .B(_03654_),
    .C(_03655_),
    .Y(_02959_)
  );
  OAI21X1 _09803_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03651_),
    .C( dbg_0.fe_mdb_in_5_ ),
    .Y(_03656_)
  );
  NOR2X1 _09804_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B( dbg_0.fe_mdb_in_4_ ),
    .Y(_03657_)
  );
  NAND2X1 _09805_ (
    .A(_03301_),
    .B(_03657_),
    .Y(_03658_)
  );
  NAND3X1 _09806_ (
    .A(_03301_),
    .B(_03644_),
    .C(_03657_),
    .Y(_03659_)
  );
  AND2X1 _09807_ (
    .A(_03656_),
    .B(_03659_),
    .Y(_03660_)
  );
  NAND2X1 _09808_ (
    .A( execution_unit_0.inst_dext_5_ ),
    .B(_03368_),
    .Y(_03661_)
  );
  OAI21X1 _09809_ (
    .A(_03368_),
    .B(_03660_),
    .C(_03661_),
    .Y(_02960_)
  );
  OR2X1 _09810_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03659_),
    .Y(_03662_)
  );
  XOR2X1 _09811_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03659_),
    .Y(_03663_)
  );
  NAND2X1 _09812_ (
    .A( execution_unit_0.inst_dext_6_ ),
    .B(_03368_),
    .Y(_03664_)
  );
  OAI21X1 _09813_ (
    .A(_03368_),
    .B(_03663_),
    .C(_03664_),
    .Y(_02961_)
  );
  NOR2X1 _09814_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03662_),
    .Y(_03665_)
  );
  XNOR2X1 _09815_ (
    .A(_03195_),
    .B(_03662_),
    .Y(_03666_)
  );
  NAND2X1 _09816_ (
    .A( execution_unit_0.inst_dext_7_ ),
    .B(_03368_),
    .Y(_03667_)
  );
  OAI21X1 _09817_ (
    .A(_03368_),
    .B(_03666_),
    .C(_03667_),
    .Y(_02962_)
  );
  OAI21X1 _09818_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03662_),
    .C( dbg_0.fe_mdb_in_8_ ),
    .Y(_03668_)
  );
  NAND2X1 _09819_ (
    .A(_03190_),
    .B(_03665_),
    .Y(_03669_)
  );
  AND2X1 _09820_ (
    .A(_03668_),
    .B(_03669_),
    .Y(_03670_)
  );
  NAND2X1 _09821_ (
    .A( execution_unit_0.inst_dext_8_ ),
    .B(_03368_),
    .Y(_03671_)
  );
  OAI21X1 _09822_ (
    .A(_03368_),
    .B(_03670_),
    .C(_03671_),
    .Y(_02963_)
  );
  NAND3X1 _09823_ (
    .A(_03190_),
    .B(_03192_),
    .C(_03195_),
    .Y(_03672_)
  );
  XNOR2X1 _09824_ (
    .A(_03192_),
    .B(_03669_),
    .Y(_03673_)
  );
  NAND2X1 _09825_ (
    .A( execution_unit_0.inst_dext_9_ ),
    .B(_03368_),
    .Y(_03674_)
  );
  OAI21X1 _09826_ (
    .A(_03368_),
    .B(_03673_),
    .C(_03674_),
    .Y(_02964_)
  );
  NOR2X1 _09827_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B( dbg_0.fe_mdb_in_6_ ),
    .Y(_03675_)
  );
  NAND3X1 _09828_ (
    .A(_03190_),
    .B(_03195_),
    .C(_03675_),
    .Y(_03676_)
  );
  NOR2X1 _09829_ (
    .A(_03658_),
    .B(_03676_),
    .Y(_03677_)
  );
  NAND2X1 _09830_ (
    .A(_03643_),
    .B(_03677_),
    .Y(_03678_)
  );
  NOR2X1 _09831_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03678_),
    .Y(_03679_)
  );
  OAI21X1 _09832_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03678_),
    .C( dbg_0.fe_mdb_in_10_ ),
    .Y(_03680_)
  );
  OR2X1 _09833_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B( dbg_0.fe_mdb_in_9_ ),
    .Y(_03681_)
  );
  OR2X1 _09834_ (
    .A(_03678_),
    .B(_03681_),
    .Y(_03682_)
  );
  AND2X1 _09835_ (
    .A(_03680_),
    .B(_03682_),
    .Y(_03683_)
  );
  NAND2X1 _09836_ (
    .A( execution_unit_0.inst_dext_10_ ),
    .B(_03368_),
    .Y(_03684_)
  );
  OAI21X1 _09837_ (
    .A(_03368_),
    .B(_03683_),
    .C(_03684_),
    .Y(_02965_)
  );
  NAND2X1 _09838_ (
    .A(_03303_),
    .B(_03679_),
    .Y(_03685_)
  );
  AOI22X1 _09839_ (
    .A(_03303_),
    .B(_03679_),
    .C(_03682_),
    .D( dbg_0.fe_mdb_in_11_ ),
    .Y(_03686_)
  );
  NAND2X1 _09840_ (
    .A( execution_unit_0.inst_dext_11_ ),
    .B(_03368_),
    .Y(_03687_)
  );
  OAI21X1 _09841_ (
    .A(_03368_),
    .B(_03686_),
    .C(_03687_),
    .Y(_02966_)
  );
  NAND2X1 _09842_ (
    .A( execution_unit_0.inst_dext_12_ ),
    .B(_03368_),
    .Y(_03688_)
  );
  OR2X1 _09843_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B( dbg_0.fe_mdb_in_12_ ),
    .Y(_03689_)
  );
  NOR2X1 _09844_ (
    .A(_03681_),
    .B(_03689_),
    .Y(_03690_)
  );
  NAND3X1 _09845_ (
    .A(_03643_),
    .B(_03677_),
    .C(_03690_),
    .Y(_03691_)
  );
  INVX1 _09846_ (
    .A(_03691_),
    .Y(_03692_)
  );
  AOI21X1 _09847_ (
    .A( dbg_0.fe_mdb_in_12_ ),
    .B(_03685_),
    .C(_03692_),
    .Y(_03693_)
  );
  OAI21X1 _09848_ (
    .A(_03368_),
    .B(_03693_),
    .C(_03688_),
    .Y(_02967_)
  );
  NAND2X1 _09849_ (
    .A( execution_unit_0.inst_dext_13_ ),
    .B(_03368_),
    .Y(_03694_)
  );
  NAND2X1 _09850_ (
    .A(_03186_),
    .B(_03692_),
    .Y(_03695_)
  );
  XNOR2X1 _09851_ (
    .A(_03186_),
    .B(_03691_),
    .Y(_03696_)
  );
  OAI21X1 _09852_ (
    .A(_03368_),
    .B(_03696_),
    .C(_03694_),
    .Y(_02968_)
  );
  AOI21X1 _09853_ (
    .A(_03186_),
    .B(_03692_),
    .C(_03185_),
    .Y(_03697_)
  );
  NOR2X1 _09854_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_03695_),
    .Y(_03698_)
  );
  OR2X1 _09855_ (
    .A(_03697_),
    .B(_03698_),
    .Y(_03699_)
  );
  OAI21X1 _09856_ (
    .A(_03697_),
    .B(_03698_),
    .C(_03369_),
    .Y(_03700_)
  );
  OAI21X1 _09857_ (
    .A(_03234_),
    .B(_03369_),
    .C(_03700_),
    .Y(_02969_)
  );
  XNOR2X1 _09858_ (
    .A(_03187_),
    .B(_03698_),
    .Y(_03701_)
  );
  NOR2X1 _09859_ (
    .A( execution_unit_0.inst_dext_15_ ),
    .B(_03369_),
    .Y(_03702_)
  );
  NOR2X1 _09860_ (
    .A(_03368_),
    .B(_03701_),
    .Y(_03703_)
  );
  NOR2X1 _09861_ (
    .A(_03702_),
    .B(_03703_),
    .Y(_02970_)
  );
  NOR2X1 _09862_ (
    .A(_03294_),
    .B(_03337_),
    .Y(_03704_)
  );
  OR2X1 _09863_ (
    .A(_03308_),
    .B(_03311_),
    .Y(_03705_)
  );
  NOR2X1 _09864_ (
    .A(_03296_),
    .B(_03705_),
    .Y(_03706_)
  );
  OAI21X1 _09865_ (
    .A(_03704_),
    .B(_03706_),
    .C(_03639_),
    .Y(_03707_)
  );
  INVX1 _09866_ (
    .A(_03707_),
    .Y(_03708_)
  );
  NOR2X1 _09867_ (
    .A(_03295_),
    .B(_03418_),
    .Y(_03709_)
  );
  OAI21X1 _09868_ (
    .A(_03295_),
    .B(_03418_),
    .C(_03374_),
    .Y(_03710_)
  );
  NOR2X1 _09869_ (
    .A(_03708_),
    .B(_03710_),
    .Y(_03711_)
  );
  NAND3X1 _09870_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03639_),
    .C(_03704_),
    .Y(_03712_)
  );
  OAI21X1 _09871_ (
    .A(_03295_),
    .B(_03418_),
    .C( dbg_0.fe_mdb_in_0_ ),
    .Y(_03713_)
  );
  OAI21X1 _09872_ (
    .A(_03708_),
    .B(_03713_),
    .C(_03712_),
    .Y(_03714_)
  );
  MUX2X1 _09873_ (
    .A( execution_unit_0.inst_sext_0_ ),
    .B(_03714_),
    .S(_03711_),
    .Y(_03715_)
  );
  INVX1 _09874_ (
    .A(_03715_),
    .Y(_02971_)
  );
  NOR2X1 _09875_ (
    .A(_03296_),
    .B(_03337_),
    .Y(_03716_)
  );
  NAND2X1 _09876_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_03709_),
    .Y(_03717_)
  );
  OAI21X1 _09877_ (
    .A(_03646_),
    .B(_03709_),
    .C(_03717_),
    .Y(_02996_)
  );
  AOI22X1 _09878_ (
    .A(_03639_),
    .B(_03716_),
    .C(_02996_),
    .D(_03707_),
    .Y(_02997_)
  );
  NAND2X1 _09879_ (
    .A( execution_unit_0.inst_sext_1_ ),
    .B(_03711_),
    .Y(_02998_)
  );
  OAI21X1 _09880_ (
    .A(_03711_),
    .B(_02997_),
    .C(_02998_),
    .Y(_02972_)
  );
  NOR2X1 _09881_ (
    .A(_03297_),
    .B(_03337_),
    .Y(_02999_)
  );
  AOI21X1 _09882_ (
    .A(_03708_),
    .B(_02999_),
    .C(_03711_),
    .Y(_03000_)
  );
  NAND2X1 _09883_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B(_03709_),
    .Y(_03001_)
  );
  OAI21X1 _09884_ (
    .A(_03648_),
    .B(_03709_),
    .C(_03001_),
    .Y(_03002_)
  );
  OAI21X1 _09885_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03323_),
    .Y(_03003_)
  );
  NOR2X1 _09886_ (
    .A(_03705_),
    .B(_03003_),
    .Y(_03004_)
  );
  AOI21X1 _09887_ (
    .A(_03707_),
    .B(_03002_),
    .C(_03004_),
    .Y(_03005_)
  );
  AOI22X1 _09888_ (
    .A(_03235_),
    .B(_03711_),
    .C(_03000_),
    .D(_03005_),
    .Y(_02973_)
  );
  OAI21X1 _09889_ (
    .A(_03297_),
    .B(_03311_),
    .C(_03708_),
    .Y(_03006_)
  );
  MUX2X1 _09890_ (
    .A(_03188_),
    .B(_03652_),
    .S(_03709_),
    .Y(_03007_)
  );
  OAI21X1 _09891_ (
    .A(_03708_),
    .B(_03007_),
    .C(_03006_),
    .Y(_03008_)
  );
  NAND2X1 _09892_ (
    .A( execution_unit_0.inst_sext_3_ ),
    .B(_03711_),
    .Y(_03009_)
  );
  OAI21X1 _09893_ (
    .A(_03711_),
    .B(_03008_),
    .C(_03009_),
    .Y(_02974_)
  );
  NAND2X1 _09894_ (
    .A( dbg_0.fe_mdb_in_3_ ),
    .B(_03709_),
    .Y(_03010_)
  );
  OAI21X1 _09895_ (
    .A(_03654_),
    .B(_03709_),
    .C(_03010_),
    .Y(_03011_)
  );
  NAND2X1 _09896_ (
    .A(_03707_),
    .B(_03011_),
    .Y(_03012_)
  );
  AOI22X1 _09897_ (
    .A(_03236_),
    .B(_03711_),
    .C(_03000_),
    .D(_03012_),
    .Y(_02975_)
  );
  NAND2X1 _09898_ (
    .A( dbg_0.fe_mdb_in_4_ ),
    .B(_03709_),
    .Y(_03013_)
  );
  OAI21X1 _09899_ (
    .A(_03660_),
    .B(_03709_),
    .C(_03013_),
    .Y(_03014_)
  );
  NAND2X1 _09900_ (
    .A(_03707_),
    .B(_03014_),
    .Y(_03015_)
  );
  AOI22X1 _09901_ (
    .A(_03237_),
    .B(_03711_),
    .C(_03000_),
    .D(_03015_),
    .Y(_02976_)
  );
  NAND2X1 _09902_ (
    .A( dbg_0.fe_mdb_in_5_ ),
    .B(_03709_),
    .Y(_03016_)
  );
  OAI21X1 _09903_ (
    .A(_03663_),
    .B(_03709_),
    .C(_03016_),
    .Y(_03017_)
  );
  NAND2X1 _09904_ (
    .A(_03707_),
    .B(_03017_),
    .Y(_03018_)
  );
  AOI22X1 _09905_ (
    .A(_03238_),
    .B(_03711_),
    .C(_03000_),
    .D(_03018_),
    .Y(_02977_)
  );
  NAND2X1 _09906_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03709_),
    .Y(_03019_)
  );
  OAI21X1 _09907_ (
    .A(_03666_),
    .B(_03709_),
    .C(_03019_),
    .Y(_03020_)
  );
  NAND2X1 _09908_ (
    .A(_03707_),
    .B(_03020_),
    .Y(_03021_)
  );
  AOI22X1 _09909_ (
    .A(_03239_),
    .B(_03711_),
    .C(_03000_),
    .D(_03021_),
    .Y(_02978_)
  );
  NAND2X1 _09910_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03709_),
    .Y(_03022_)
  );
  OAI21X1 _09911_ (
    .A(_03670_),
    .B(_03709_),
    .C(_03022_),
    .Y(_03023_)
  );
  NAND2X1 _09912_ (
    .A(_03707_),
    .B(_03023_),
    .Y(_03024_)
  );
  AOI22X1 _09913_ (
    .A(_03240_),
    .B(_03711_),
    .C(_03000_),
    .D(_03024_),
    .Y(_02979_)
  );
  NAND2X1 _09914_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03709_),
    .Y(_03025_)
  );
  OAI21X1 _09915_ (
    .A(_03673_),
    .B(_03709_),
    .C(_03025_),
    .Y(_03026_)
  );
  NAND2X1 _09916_ (
    .A(_03707_),
    .B(_03026_),
    .Y(_03027_)
  );
  AOI22X1 _09917_ (
    .A(_03241_),
    .B(_03711_),
    .C(_03000_),
    .D(_03027_),
    .Y(_02980_)
  );
  NOR2X1 _09918_ (
    .A(_03683_),
    .B(_03709_),
    .Y(_03028_)
  );
  AND2X1 _09919_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03709_),
    .Y(_03029_)
  );
  OAI21X1 _09920_ (
    .A(_03028_),
    .B(_03029_),
    .C(_03707_),
    .Y(_03030_)
  );
  AOI22X1 _09921_ (
    .A(_03242_),
    .B(_03711_),
    .C(_03000_),
    .D(_03030_),
    .Y(_02981_)
  );
  NOR2X1 _09922_ (
    .A(_03686_),
    .B(_03709_),
    .Y(_03031_)
  );
  OAI21X1 _09923_ (
    .A(_03029_),
    .B(_03031_),
    .C(_03707_),
    .Y(_03032_)
  );
  AOI22X1 _09924_ (
    .A(_03243_),
    .B(_03711_),
    .C(_03000_),
    .D(_03032_),
    .Y(_02982_)
  );
  NOR2X1 _09925_ (
    .A(_03693_),
    .B(_03709_),
    .Y(_03033_)
  );
  OAI21X1 _09926_ (
    .A(_03029_),
    .B(_03033_),
    .C(_03707_),
    .Y(_03034_)
  );
  AOI22X1 _09927_ (
    .A(_03244_),
    .B(_03711_),
    .C(_03000_),
    .D(_03034_),
    .Y(_02983_)
  );
  NOR2X1 _09928_ (
    .A(_03696_),
    .B(_03709_),
    .Y(_03035_)
  );
  OAI21X1 _09929_ (
    .A(_03029_),
    .B(_03035_),
    .C(_03707_),
    .Y(_03036_)
  );
  AOI22X1 _09930_ (
    .A(_03245_),
    .B(_03711_),
    .C(_03000_),
    .D(_03036_),
    .Y(_02984_)
  );
  OAI21X1 _09931_ (
    .A(_03699_),
    .B(_03029_),
    .C(_03707_),
    .Y(_03037_)
  );
  AOI22X1 _09932_ (
    .A(_03246_),
    .B(_03711_),
    .C(_03000_),
    .D(_03037_),
    .Y(_02985_)
  );
  OAI21X1 _09933_ (
    .A(_03701_),
    .B(_03029_),
    .C(_03707_),
    .Y(_03038_)
  );
  AOI22X1 _09934_ (
    .A(_03247_),
    .B(_03711_),
    .C(_03000_),
    .D(_03038_),
    .Y(_02986_)
  );
  AND2X1 _09935_ (
    .A( execution_unit_0.inst_irq_rst ),
    .B(_03268_),
    .Y(_02991_)
  );
  NOR2X1 _09936_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B( dbg_0.fe_mdb_in_12_ ),
    .Y(_03039_)
  );
  INVX1 _09937_ (
    .A(_03039_),
    .Y(_03040_)
  );
  NAND2X1 _09938_ (
    .A( dbg_0.fe_mdb_in_15_ ),
    .B(_03291_),
    .Y(_03041_)
  );
  INVX1 _09939_ (
    .A(_03041_),
    .Y(_03042_)
  );
  NAND2X1 _09940_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_03042_),
    .Y(_03043_)
  );
  NOR2X1 _09941_ (
    .A(_03040_),
    .B(_03043_),
    .Y(_03044_)
  );
  NAND2X1 _09942_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B( dbg_0.fe_mdb_in_12_ ),
    .Y(_03045_)
  );
  NAND2X1 _09943_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B(_03187_),
    .Y(_03046_)
  );
  NOR2X1 _09944_ (
    .A( dbg_0.fe_mdb_in_13_ ),
    .B(_03187_),
    .Y(_03047_)
  );
  NAND2X1 _09945_ (
    .A(_03185_),
    .B(_03047_),
    .Y(_03048_)
  );
  OAI21X1 _09946_ (
    .A(_03045_),
    .B(_03046_),
    .C(_03048_),
    .Y(_03049_)
  );
  AOI21X1 _09947_ (
    .A(_03291_),
    .B(_03049_),
    .C(_03044_),
    .Y(_03050_)
  );
  NAND2X1 _09948_ (
    .A( execution_unit_0.alu_0.inst_alu_0_ ),
    .B(_03638_),
    .Y(_03051_)
  );
  OAI21X1 _09949_ (
    .A(_03638_),
    .B(_03050_),
    .C(_03051_),
    .Y(_02908_)
  );
  NAND2X1 _09950_ (
    .A( execution_unit_0.alu_0.inst_alu_1_ ),
    .B(_03638_),
    .Y(_03052_)
  );
  OAI21X1 _09951_ (
    .A(_03421_),
    .B(_03048_),
    .C(_03052_),
    .Y(_02909_)
  );
  NOR2X1 _09952_ (
    .A(_03186_),
    .B(_03046_),
    .Y(_03053_)
  );
  AOI22X1 _09953_ (
    .A( execution_unit_0.alu_0.inst_alu_2_ ),
    .B(_03638_),
    .C(_03053_),
    .D(_03420_),
    .Y(_03054_)
  );
  NAND2X1 _09954_ (
    .A(_03185_),
    .B(_03042_),
    .Y(_03055_)
  );
  NOR2X1 _09955_ (
    .A(_03186_),
    .B( dbg_0.fe_mdb_in_12_ ),
    .Y(_03056_)
  );
  NAND2X1 _09956_ (
    .A( dbg_0.decode_noirq ),
    .B(_03056_),
    .Y(_03057_)
  );
  OAI21X1 _09957_ (
    .A(_03055_),
    .B(_03057_),
    .C(_03054_),
    .Y(_02910_)
  );
  OAI21X1 _09958_ (
    .A(_03039_),
    .B(_03046_),
    .C(_03048_),
    .Y(_03058_)
  );
  OAI21X1 _09959_ (
    .A(_03418_),
    .B(_03058_),
    .C(_03291_),
    .Y(_03059_)
  );
  NOR2X1 _09960_ (
    .A( execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_03639_),
    .Y(_03060_)
  );
  AOI21X1 _09961_ (
    .A(_03633_),
    .B(_03059_),
    .C(_03060_),
    .Y(_02911_)
  );
  NOR2X1 _09962_ (
    .A(_03041_),
    .B(_03045_),
    .Y(_03061_)
  );
  OAI21X1 _09963_ (
    .A(_03044_),
    .B(_03061_),
    .C(_03639_),
    .Y(_03062_)
  );
  OAI21X1 _09964_ (
    .A(_03248_),
    .B(_03639_),
    .C(_03062_),
    .Y(_02912_)
  );
  NAND2X1 _09965_ (
    .A( execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_03638_),
    .Y(_03063_)
  );
  OAI21X1 _09966_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.fe_mdb_in_15_ ),
    .C(_03420_),
    .Y(_03064_)
  );
  NAND3X1 _09967_ (
    .A( dbg_0.fe_mdb_in_14_ ),
    .B( dbg_0.fe_mdb_in_12_ ),
    .C(_03047_),
    .Y(_03065_)
  );
  OAI21X1 _09968_ (
    .A(_03064_),
    .B(_03065_),
    .C(_03063_),
    .Y(_02913_)
  );
  NAND2X1 _09969_ (
    .A( execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_03638_),
    .Y(_03066_)
  );
  OAI21X1 _09970_ (
    .A(_03043_),
    .B(_03057_),
    .C(_03066_),
    .Y(_02914_)
  );
  NAND2X1 _09971_ (
    .A( execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_03638_),
    .Y(_03067_)
  );
  OAI21X1 _09972_ (
    .A(_03055_),
    .B(_03057_),
    .C(_03067_),
    .Y(_02915_)
  );
  AOI22X1 _09973_ (
    .A( execution_unit_0.alu_0.inst_alu_8_ ),
    .B(_03638_),
    .C(_03061_),
    .D( dbg_0.decode_noirq ),
    .Y(_03068_)
  );
  NOR2X1 _09974_ (
    .A( dbg_0.fe_mdb_in_9_ ),
    .B(_03638_),
    .Y(_03069_)
  );
  NAND2X1 _09975_ (
    .A(_03300_),
    .B(_03069_),
    .Y(_03070_)
  );
  OAI21X1 _09976_ (
    .A(_03352_),
    .B(_03070_),
    .C(_03068_),
    .Y(_02916_)
  );
  OAI21X1 _09977_ (
    .A( dbg_0.fe_mdb_in_8_ ),
    .B(_03195_),
    .C(_03192_),
    .Y(_03071_)
  );
  NOR2X1 _09978_ (
    .A(_03299_),
    .B(_03071_),
    .Y(_03072_)
  );
  OAI21X1 _09979_ (
    .A(_03186_),
    .B(_03041_),
    .C(_03059_),
    .Y(_03073_)
  );
  OAI22X1 _09980_ (
    .A( execution_unit_0.alu_0.inst_alu_9_ ),
    .B(_03639_),
    .C(_03072_),
    .D(_03073_),
    .Y(_03074_)
  );
  INVX1 _09981_ (
    .A(_03074_),
    .Y(_02917_)
  );
  NAND2X1 _09982_ (
    .A( execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_03638_),
    .Y(_03075_)
  );
  OAI21X1 _09983_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03070_),
    .C(_03075_),
    .Y(_02918_)
  );
  OAI21X1 _09984_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C( dbg_0.fe_mdb_in_12_ ),
    .Y(_03076_)
  );
  NAND2X1 _09985_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_03638_),
    .Y(_03077_)
  );
  OAI21X1 _09986_ (
    .A(_03055_),
    .B(_03076_),
    .C(_03077_),
    .Y(_02919_)
  );
  OAI21X1 _09987_ (
    .A(_03331_),
    .B(_03388_),
    .C(_03639_),
    .Y(_03078_)
  );
  NAND2X1 _09988_ (
    .A( frontend_0.inst_sz_0_ ),
    .B(_03638_),
    .Y(_03079_)
  );
  OAI21X1 _09989_ (
    .A(_03414_),
    .B(_03078_),
    .C(_03079_),
    .Y(_02924_)
  );
  OAI21X1 _09990_ (
    .A( frontend_0.inst_sz_1_ ),
    .B(_03639_),
    .C(_03078_),
    .Y(_03080_)
  );
  INVX1 _09991_ (
    .A(_03080_),
    .Y(_02925_)
  );
  NAND2X1 _09992_ (
    .A( dbg_0.fe_mdb_in_6_ ),
    .B(_03420_),
    .Y(_03081_)
  );
  NOR2X1 _09993_ (
    .A(_03286_),
    .B(_03081_),
    .Y(_03082_)
  );
  AOI22X1 _09994_ (
    .A( execution_unit_0.alu_0.inst_bw ),
    .B(_03638_),
    .C(_03082_),
    .D(_03295_),
    .Y(_03083_)
  );
  INVX1 _09995_ (
    .A(_03083_),
    .Y(_02926_)
  );
  AOI21X1 _09996_ (
    .A(_03337_),
    .B(_03657_),
    .C(_03294_),
    .Y(_03084_)
  );
  NAND2X1 _09997_ (
    .A( execution_unit_0.inst_as_0_ ),
    .B(_03638_),
    .Y(_03085_)
  );
  OAI21X1 _09998_ (
    .A(_03638_),
    .B(_03084_),
    .C(_03085_),
    .Y(_02927_)
  );
  OAI21X1 _09999_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03339_),
    .Y(_03086_)
  );
  NAND2X1 _10000_ (
    .A( execution_unit_0.inst_as_1_ ),
    .B(_03638_),
    .Y(_03087_)
  );
  OAI21X1 _10001_ (
    .A(_03312_),
    .B(_03086_),
    .C(_03087_),
    .Y(_02928_)
  );
  NAND2X1 _10002_ (
    .A( execution_unit_0.inst_as_2_ ),
    .B(_03638_),
    .Y(_03088_)
  );
  OAI21X1 _10003_ (
    .A(_03324_),
    .B(_03638_),
    .C(_03088_),
    .Y(_02929_)
  );
  NAND2X1 _10004_ (
    .A( execution_unit_0.inst_as_3_ ),
    .B(_03638_),
    .Y(_03089_)
  );
  OAI21X1 _10005_ (
    .A(_03314_),
    .B(_03638_),
    .C(_03089_),
    .Y(_02930_)
  );
  OAI22X1 _10006_ (
    .A(_03196_),
    .B(_03639_),
    .C(_03086_),
    .D(_03316_),
    .Y(_02931_)
  );
  NAND2X1 _10007_ (
    .A( execution_unit_0.inst_as_5_ ),
    .B(_03638_),
    .Y(_03090_)
  );
  OAI21X1 _10008_ (
    .A(_03318_),
    .B(_03638_),
    .C(_03090_),
    .Y(_02932_)
  );
  NAND2X1 _10009_ (
    .A( execution_unit_0.inst_as_6_ ),
    .B(_03638_),
    .Y(_03091_)
  );
  OAI21X1 _10010_ (
    .A(_03705_),
    .B(_03086_),
    .C(_03091_),
    .Y(_02933_)
  );
  OAI21X1 _10011_ (
    .A(_03249_),
    .B(_03639_),
    .C(_03707_),
    .Y(_02934_)
  );
  OAI21X1 _10012_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03190_),
    .Y(_03092_)
  );
  OAI21X1 _10013_ (
    .A( frontend_0.inst_src_bin_0_ ),
    .B(_03639_),
    .C(_03092_),
    .Y(_03093_)
  );
  INVX1 _10014_ (
    .A(_03093_),
    .Y(_02935_)
  );
  AOI21X1 _10015_ (
    .A(_03229_),
    .B(_03638_),
    .C(_03069_),
    .Y(_02936_)
  );
  OAI21X1 _10016_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03191_),
    .Y(_03094_)
  );
  OAI21X1 _10017_ (
    .A( frontend_0.inst_dest_bin_0_ ),
    .B(_03639_),
    .C(_03094_),
    .Y(_03095_)
  );
  INVX1 _10018_ (
    .A(_03095_),
    .Y(_02937_)
  );
  OAI21X1 _10019_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03193_),
    .Y(_03096_)
  );
  OAI21X1 _10020_ (
    .A( frontend_0.inst_dest_bin_1_ ),
    .B(_03639_),
    .C(_03096_),
    .Y(_03097_)
  );
  INVX1 _10021_ (
    .A(_03097_),
    .Y(_02938_)
  );
  OAI21X1 _10022_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03188_),
    .Y(_03098_)
  );
  OAI21X1 _10023_ (
    .A( frontend_0.inst_dest_bin_2_ ),
    .B(_03639_),
    .C(_03098_),
    .Y(_03099_)
  );
  INVX1 _10024_ (
    .A(_03099_),
    .Y(_02939_)
  );
  OAI21X1 _10025_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C(_03189_),
    .Y(_03100_)
  );
  OAI21X1 _10026_ (
    .A( frontend_0.inst_dest_bin_3_ ),
    .B(_03639_),
    .C(_03100_),
    .Y(_03101_)
  );
  INVX1 _10027_ (
    .A(_03101_),
    .Y(_02940_)
  );
  NAND2X1 _10028_ (
    .A( execution_unit_0.inst_mov ),
    .B(_03638_),
    .Y(_03102_)
  );
  NAND2X1 _10029_ (
    .A(_03420_),
    .B(_03039_),
    .Y(_03103_)
  );
  OAI21X1 _10030_ (
    .A(_03046_),
    .B(_03103_),
    .C(_03102_),
    .Y(_02941_)
  );
  MUX2X1 _10031_ (
    .A( dbg_0.fe_mdb_in_10_ ),
    .B( frontend_0.inst_jmp_bin_0_ ),
    .S(_03639_),
    .Y(_03104_)
  );
  INVX1 _10032_ (
    .A(_03104_),
    .Y(_02942_)
  );
  MUX2X1 _10033_ (
    .A( dbg_0.fe_mdb_in_11_ ),
    .B( frontend_0.inst_jmp_bin_1_ ),
    .S(_03639_),
    .Y(_03105_)
  );
  INVX1 _10034_ (
    .A(_03105_),
    .Y(_02943_)
  );
  OAI21X1 _10035_ (
    .A(_03233_),
    .B(_03639_),
    .C(_03076_),
    .Y(_02944_)
  );
  NAND2X1 _10036_ (
    .A( execution_unit_0.alu_0.inst_so_0_ ),
    .B(_03638_),
    .Y(_03106_)
  );
  NAND2X1 _10037_ (
    .A(_03300_),
    .B( dbg_0.decode_noirq ),
    .Y(_03107_)
  );
  OAI21X1 _10038_ (
    .A(_03672_),
    .B(_03107_),
    .C(_03106_),
    .Y(_02945_)
  );
  NAND2X1 _10039_ (
    .A( execution_unit_0.alu_0.inst_so_1_ ),
    .B(_03638_),
    .Y(_03108_)
  );
  NAND3X1 _10040_ (
    .A(_03190_),
    .B(_03192_),
    .C( dbg_0.fe_mdb_in_7_ ),
    .Y(_03109_)
  );
  OAI21X1 _10041_ (
    .A(_03107_),
    .B(_03109_),
    .C(_03108_),
    .Y(_02946_)
  );
  NAND2X1 _10042_ (
    .A( execution_unit_0.alu_0.inst_so_3_ ),
    .B(_03638_),
    .Y(_03110_)
  );
  OAI21X1 _10043_ (
    .A(_03352_),
    .B(_03070_),
    .C(_03110_),
    .Y(_02947_)
  );
  NAND2X1 _10044_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B(_03638_),
    .Y(_03111_)
  );
  NAND3X1 _10045_ (
    .A(_03190_),
    .B(_03320_),
    .C(_03639_),
    .Y(_03112_)
  );
  OAI21X1 _10046_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03112_),
    .C(_03111_),
    .Y(_02948_)
  );
  NAND2X1 _10047_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_03638_),
    .Y(_03113_)
  );
  OAI21X1 _10048_ (
    .A(_03195_),
    .B(_03112_),
    .C(_03113_),
    .Y(_02949_)
  );
  NAND2X1 _10049_ (
    .A( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_03638_),
    .Y(_03114_)
  );
  OAI21X1 _10050_ (
    .A(_03322_),
    .B(_03638_),
    .C(_03114_),
    .Y(_02950_)
  );
  AOI22X1 _10051_ (
    .A(_03353_),
    .B(_03420_),
    .C(_03638_),
    .D(_03223_),
    .Y(_02951_)
  );
  OAI21X1 _10052_ (
    .A(_03201_),
    .B(_03639_),
    .C(_03107_),
    .Y(_02952_)
  );
  AOI21X1 _10053_ (
    .A( execution_unit_0.inst_type_1_ ),
    .B(_03638_),
    .C(_03709_),
    .Y(_03115_)
  );
  INVX1 _10054_ (
    .A(_03115_),
    .Y(_02953_)
  );
  OAI21X1 _10055_ (
    .A(_03231_),
    .B(_03639_),
    .C(_03064_),
    .Y(_02954_)
  );
  NAND2X1 _10056_ (
    .A( execution_unit_0.inst_ad_0_ ),
    .B(_03638_),
    .Y(_03116_)
  );
  OAI21X1 _10057_ (
    .A( dbg_0.fe_mdb_in_7_ ),
    .B(_03064_),
    .C(_03116_),
    .Y(_02987_)
  );
  OAI21X1 _10058_ (
    .A(_03290_),
    .B( dbg_0.decode_noirq ),
    .C( dbg_0.fe_mdb_in_7_ ),
    .Y(_03117_)
  );
  OAI21X1 _10059_ (
    .A( dbg_0.fe_mdb_in_0_ ),
    .B(_03302_),
    .C(_03329_),
    .Y(_03118_)
  );
  OAI22X1 _10060_ (
    .A(_03198_),
    .B(_03639_),
    .C(_03117_),
    .D(_03118_),
    .Y(_02988_)
  );
  NAND2X1 _10061_ (
    .A( execution_unit_0.UNUSED_inst_ad_symb ),
    .B(_03638_),
    .Y(_03119_)
  );
  OAI21X1 _10062_ (
    .A(_03635_),
    .B(_03117_),
    .C(_03119_),
    .Y(_02989_)
  );
  NAND2X1 _10063_ (
    .A( execution_unit_0.inst_ad_6_ ),
    .B(_03638_),
    .Y(_03120_)
  );
  NAND3X1 _10064_ (
    .A( dbg_0.fe_mdb_in_1_ ),
    .B(_03301_),
    .C(_03330_),
    .Y(_03121_)
  );
  OAI21X1 _10065_ (
    .A(_03094_),
    .B(_03121_),
    .C(_03120_),
    .Y(_02990_)
  );
  NOR2X1 _10066_ (
    .A(1'h0),
    .B(_03281_),
    .Y(_03122_)
  );
  NAND3X1 _10067_ (
    .A(_03173_),
    .B(irq_8_),
    .C(_03273_),
    .Y(_03123_)
  );
  OAI21X1 _10068_ (
    .A(irq_10_),
    .B( frontend_0.wdt_irq ),
    .C(_03174_),
    .Y(_03124_)
  );
  AOI21X1 _10069_ (
    .A(_03175_),
    .B(_03124_),
    .C(irq_13_),
    .Y(_03125_)
  );
  OAI21X1 _10070_ (
    .A(_03281_),
    .B(_03123_),
    .C(_03177_),
    .Y(_03126_)
  );
  NOR2X1 _10071_ (
    .A(_03125_),
    .B(_03126_),
    .Y(_03127_)
  );
  AND2X1 _10072_ (
    .A(_03275_),
    .B(_03122_),
    .Y(_03128_)
  );
  OAI21X1 _10073_ (
    .A(irq_9_),
    .B(irq_8_),
    .C(_03273_),
    .Y(_03129_)
  );
  AOI21X1 _10074_ (
    .A(_03280_),
    .B(_03129_),
    .C(1'h0),
    .Y(_03130_)
  );
  INVX1 _10075_ (
    .A(_03130_),
    .Y(_03131_)
  );
  NOR2X1 _10076_ (
    .A(_03128_),
    .B(_03130_),
    .Y(_03132_)
  );
  NAND3X1 _10077_ (
    .A(_03172_),
    .B(irq_6_),
    .C(_03132_),
    .Y(_03133_)
  );
  AND2X1 _10078_ (
    .A(_03127_),
    .B(_03133_),
    .Y(_03134_)
  );
  NAND2X1 _10079_ (
    .A(_03171_),
    .B(_03279_),
    .Y(_03135_)
  );
  AND2X1 _10080_ (
    .A(_03127_),
    .B(_03132_),
    .Y(_03136_)
  );
  NAND2X1 _10081_ (
    .A(irq_4_),
    .B(_03136_),
    .Y(_03137_)
  );
  NOR2X1 _10082_ (
    .A(_03135_),
    .B(_03137_),
    .Y(_03138_)
  );
  OAI21X1 _10083_ (
    .A(_03135_),
    .B(_03137_),
    .C(_03134_),
    .Y(_03139_)
  );
  INVX1 _10084_ (
    .A(_03139_),
    .Y(_03140_)
  );
  OAI21X1 _10085_ (
    .A(irq_4_),
    .B(_03135_),
    .C(_03136_),
    .Y(_03141_)
  );
  NAND2X1 _10086_ (
    .A(_03132_),
    .B(_03141_),
    .Y(_03142_)
  );
  NOR2X1 _10087_ (
    .A(_03139_),
    .B(_03142_),
    .Y(_03143_)
  );
  NAND2X1 _10088_ (
    .A(irq_2_),
    .B(_03143_),
    .Y(_03144_)
  );
  OAI21X1 _10089_ (
    .A(irq_3_),
    .B(irq_2_),
    .C(_03143_),
    .Y(_03145_)
  );
  INVX1 _10090_ (
    .A(_03145_),
    .Y(_03146_)
  );
  NAND2X1 _10091_ (
    .A(_03141_),
    .B(_03145_),
    .Y(_03147_)
  );
  OAI21X1 _10092_ (
    .A(irq_3_),
    .B(_03144_),
    .C(_03140_),
    .Y(_03148_)
  );
  OR2X1 _10093_ (
    .A(_03139_),
    .B(_03147_),
    .Y(_03149_)
  );
  INVX1 _10094_ (
    .A(_03149_),
    .Y(_03150_)
  );
  NOR2X1 _10095_ (
    .A(_03128_),
    .B(_03146_),
    .Y(_03151_)
  );
  INVX1 _10096_ (
    .A(_03151_),
    .Y(_03152_)
  );
  NAND3X1 _10097_ (
    .A(irq_5_),
    .B(_03279_),
    .C(_03136_),
    .Y(_03153_)
  );
  NAND2X1 _10098_ (
    .A(_03131_),
    .B(_03153_),
    .Y(_03154_)
  );
  NOR2X1 _10099_ (
    .A(_03138_),
    .B(_03154_),
    .Y(_03155_)
  );
  NAND3X1 _10100_ (
    .A(irq_1_),
    .B(_03151_),
    .C(_03155_),
    .Y(_03156_)
  );
  OR2X1 _10101_ (
    .A(_03149_),
    .B(_03156_),
    .Y(_03157_)
  );
  NAND3X1 _10102_ (
    .A(irq_0_),
    .B(_03150_),
    .C(_03151_),
    .Y(_03158_)
  );
  OAI21X1 _10103_ (
    .A(_03149_),
    .B(_03156_),
    .C(_03155_),
    .Y(_03159_)
  );
  OR2X1 _10104_ (
    .A(_03158_),
    .B(_03159_),
    .Y(_03160_)
  );
  NOR2X1 _10105_ (
    .A(_03291_),
    .B(_03148_),
    .Y(_03161_)
  );
  AOI22X1 _10106_ (
    .A( frontend_0.irq_addr_1_ ),
    .B(_03291_),
    .C(_03160_),
    .D(_03161_),
    .Y(_03162_)
  );
  INVX1 _10107_ (
    .A(_03162_),
    .Y(_02992_)
  );
  NAND2X1 _10108_ (
    .A( frontend_0.irq_addr_2_ ),
    .B(_03291_),
    .Y(_03163_)
  );
  NAND3X1 _10109_ (
    .A(_03155_),
    .B(_03157_),
    .C(_03158_),
    .Y(_03164_)
  );
  OAI21X1 _10110_ (
    .A(_03291_),
    .B(_03164_),
    .C(_03163_),
    .Y(_02993_)
  );
  NAND3X1 _10111_ (
    .A(_03290_),
    .B(_03157_),
    .C(_03160_),
    .Y(_03165_)
  );
  OAI22X1 _10112_ (
    .A(_03208_),
    .B(_03290_),
    .C(_03152_),
    .D(_03165_),
    .Y(_02994_)
  );
  NAND2X1 _10113_ (
    .A( frontend_0.irq_addr_4_ ),
    .B(_03291_),
    .Y(_03166_)
  );
  OAI21X1 _10114_ (
    .A(_03147_),
    .B(_03165_),
    .C(_03166_),
    .Y(_02995_)
  );
  DFFSR _10115_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_0_ ),
    .Q( execution_unit_0.e_state_0_ ),
    .R(1'h1),
    .S(_02907_)
  );
  DFFSR _10116_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_1_ ),
    .Q( execution_unit_0.e_state_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10117_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_2_ ),
    .Q( execution_unit_0.e_state_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10118_ (
    .CLK(dco_clk),
    .D( frontend_0.e_state_nxt_3_ ),
    .Q( execution_unit_0.e_state_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10119_ (
    .CLK(dco_clk),
    .D(_02908_),
    .Q( execution_unit_0.alu_0.inst_alu_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10120_ (
    .CLK(dco_clk),
    .D(_02909_),
    .Q( execution_unit_0.alu_0.inst_alu_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10121_ (
    .CLK(dco_clk),
    .D(_02910_),
    .Q( execution_unit_0.alu_0.inst_alu_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10122_ (
    .CLK(dco_clk),
    .D(_02911_),
    .Q( execution_unit_0.alu_0.inst_alu_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10123_ (
    .CLK(dco_clk),
    .D(_02912_),
    .Q( execution_unit_0.alu_0.inst_alu_4_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10124_ (
    .CLK(dco_clk),
    .D(_02913_),
    .Q( execution_unit_0.alu_0.inst_alu_5_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10125_ (
    .CLK(dco_clk),
    .D(_02914_),
    .Q( execution_unit_0.alu_0.inst_alu_6_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10126_ (
    .CLK(dco_clk),
    .D(_02915_),
    .Q( execution_unit_0.alu_0.inst_alu_7_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10127_ (
    .CLK(dco_clk),
    .D(_02916_),
    .Q( execution_unit_0.alu_0.inst_alu_8_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10128_ (
    .CLK(dco_clk),
    .D(_02917_),
    .Q( execution_unit_0.alu_0.inst_alu_9_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10129_ (
    .CLK(dco_clk),
    .D(_02918_),
    .Q( execution_unit_0.alu_0.inst_alu_10_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10130_ (
    .CLK(dco_clk),
    .D(_02919_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_alu ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10131_ (
    .CLK(dco_clk),
    .D(_02920_),
    .Q( frontend_0.exec_dext_rdy ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10132_ (
    .CLK(dco_clk),
    .D(_02921_),
    .Q( frontend_0.exec_src_wr ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10133_ (
    .CLK(dco_clk),
    .D(_02922_),
    .Q( frontend_0.exec_dst_wr ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10134_ (
    .CLK(dco_clk),
    .D(_02923_),
    .Q( frontend_0.exec_jmp ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10135_ (
    .CLK(dco_clk),
    .D(_02924_),
    .Q( frontend_0.inst_sz_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10136_ (
    .CLK(dco_clk),
    .D(_02925_),
    .Q( frontend_0.inst_sz_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10137_ (
    .CLK(dco_clk),
    .D(_02926_),
    .Q( execution_unit_0.alu_0.inst_bw ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10138_ (
    .CLK(dco_clk),
    .D(_02927_),
    .Q( execution_unit_0.inst_as_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10139_ (
    .CLK(dco_clk),
    .D(_02928_),
    .Q( execution_unit_0.inst_as_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10140_ (
    .CLK(dco_clk),
    .D(_02929_),
    .Q( execution_unit_0.inst_as_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10141_ (
    .CLK(dco_clk),
    .D(_02930_),
    .Q( execution_unit_0.inst_as_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10142_ (
    .CLK(dco_clk),
    .D(_02931_),
    .Q( execution_unit_0.inst_as_4_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10143_ (
    .CLK(dco_clk),
    .D(_02932_),
    .Q( execution_unit_0.inst_as_5_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10144_ (
    .CLK(dco_clk),
    .D(_02933_),
    .Q( execution_unit_0.inst_as_6_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10145_ (
    .CLK(dco_clk),
    .D(_02934_),
    .Q( execution_unit_0.inst_as_7_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10146_ (
    .CLK(dco_clk),
    .D(_02935_),
    .Q( frontend_0.inst_src_bin_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10147_ (
    .CLK(dco_clk),
    .D(_02936_),
    .Q( frontend_0.inst_src_bin_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10148_ (
    .CLK(dco_clk),
    .D(_02937_),
    .Q( frontend_0.inst_dest_bin_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10149_ (
    .CLK(dco_clk),
    .D(_02938_),
    .Q( frontend_0.inst_dest_bin_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10150_ (
    .CLK(dco_clk),
    .D(_02939_),
    .Q( frontend_0.inst_dest_bin_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10151_ (
    .CLK(dco_clk),
    .D(_02940_),
    .Q( frontend_0.inst_dest_bin_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10152_ (
    .CLK(dco_clk),
    .D(_02941_),
    .Q( execution_unit_0.inst_mov ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10153_ (
    .CLK(dco_clk),
    .D(_02942_),
    .Q( frontend_0.inst_jmp_bin_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10154_ (
    .CLK(dco_clk),
    .D(_02943_),
    .Q( frontend_0.inst_jmp_bin_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10155_ (
    .CLK(dco_clk),
    .D(_02944_),
    .Q( frontend_0.inst_jmp_bin_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10156_ (
    .CLK(dco_clk),
    .D(_02945_),
    .Q( execution_unit_0.alu_0.inst_so_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10157_ (
    .CLK(dco_clk),
    .D(_02946_),
    .Q( execution_unit_0.alu_0.inst_so_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10158_ (
    .CLK(dco_clk),
    .D(_02947_),
    .Q( execution_unit_0.alu_0.inst_so_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10159_ (
    .CLK(dco_clk),
    .D(_02948_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10160_ (
    .CLK(dco_clk),
    .D(_02949_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10161_ (
    .CLK(dco_clk),
    .D(_02950_),
    .Q( execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10162_ (
    .CLK(dco_clk),
    .D(_02951_),
    .Q( execution_unit_0.alu_0.inst_so_7_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10163_ (
    .CLK(dco_clk),
    .D(_02952_),
    .Q( execution_unit_0.inst_type_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10164_ (
    .CLK(dco_clk),
    .D(_02953_),
    .Q( execution_unit_0.inst_type_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10165_ (
    .CLK(dco_clk),
    .D(_02954_),
    .Q( execution_unit_0.inst_type_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10166_ (
    .CLK(dco_clk),
    .D(_02955_),
    .Q( execution_unit_0.inst_dext_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10167_ (
    .CLK(dco_clk),
    .D(_02956_),
    .Q( execution_unit_0.inst_dext_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10168_ (
    .CLK(dco_clk),
    .D(_02957_),
    .Q( execution_unit_0.inst_dext_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10169_ (
    .CLK(dco_clk),
    .D(_02958_),
    .Q( execution_unit_0.inst_dext_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10170_ (
    .CLK(dco_clk),
    .D(_02959_),
    .Q( execution_unit_0.inst_dext_4_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10171_ (
    .CLK(dco_clk),
    .D(_02960_),
    .Q( execution_unit_0.inst_dext_5_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10172_ (
    .CLK(dco_clk),
    .D(_02961_),
    .Q( execution_unit_0.inst_dext_6_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10173_ (
    .CLK(dco_clk),
    .D(_02962_),
    .Q( execution_unit_0.inst_dext_7_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10174_ (
    .CLK(dco_clk),
    .D(_02963_),
    .Q( execution_unit_0.inst_dext_8_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10175_ (
    .CLK(dco_clk),
    .D(_02964_),
    .Q( execution_unit_0.inst_dext_9_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10176_ (
    .CLK(dco_clk),
    .D(_02965_),
    .Q( execution_unit_0.inst_dext_10_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10177_ (
    .CLK(dco_clk),
    .D(_02966_),
    .Q( execution_unit_0.inst_dext_11_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10178_ (
    .CLK(dco_clk),
    .D(_02967_),
    .Q( execution_unit_0.inst_dext_12_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10179_ (
    .CLK(dco_clk),
    .D(_02968_),
    .Q( execution_unit_0.inst_dext_13_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10180_ (
    .CLK(dco_clk),
    .D(_02969_),
    .Q( execution_unit_0.inst_dext_14_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10181_ (
    .CLK(dco_clk),
    .D(_02970_),
    .Q( execution_unit_0.inst_dext_15_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10182_ (
    .CLK(dco_clk),
    .D( frontend_0.fe_pmem_wait ),
    .Q( frontend_0.pmem_busy ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10183_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_0_ ),
    .Q( dbg_0.UNUSED_pc_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10184_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_1_ ),
    .Q( dbg_0.UNUSED_pc_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10185_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_2_ ),
    .Q( dbg_0.UNUSED_pc_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10186_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_3_ ),
    .Q( dbg_0.UNUSED_pc_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10187_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_4_ ),
    .Q( dbg_0.UNUSED_pc_4_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10188_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_5_ ),
    .Q( dbg_0.UNUSED_pc_5_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10189_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_6_ ),
    .Q( dbg_0.UNUSED_pc_6_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10190_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_7_ ),
    .Q( dbg_0.UNUSED_pc_7_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10191_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_8_ ),
    .Q( dbg_0.UNUSED_pc_8_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10192_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_9_ ),
    .Q( dbg_0.UNUSED_pc_9_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10193_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_10_ ),
    .Q( dbg_0.UNUSED_pc_10_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10194_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_11_ ),
    .Q( dbg_0.UNUSED_pc_11_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10195_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_12_ ),
    .Q( dbg_0.UNUSED_pc_12_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10196_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_13_ ),
    .Q( dbg_0.UNUSED_pc_13_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10197_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_14_ ),
    .Q( dbg_0.UNUSED_pc_14_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10198_ (
    .CLK(dco_clk),
    .D( execution_unit_0.pc_nxt_15_ ),
    .Q( dbg_0.UNUSED_pc_15_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10199_ (
    .CLK(dco_clk),
    .D(_02971_),
    .Q( execution_unit_0.inst_sext_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10200_ (
    .CLK(dco_clk),
    .D(_02972_),
    .Q( execution_unit_0.inst_sext_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10201_ (
    .CLK(dco_clk),
    .D(_02973_),
    .Q( execution_unit_0.inst_sext_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10202_ (
    .CLK(dco_clk),
    .D(_02974_),
    .Q( execution_unit_0.inst_sext_3_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10203_ (
    .CLK(dco_clk),
    .D(_02975_),
    .Q( execution_unit_0.inst_sext_4_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10204_ (
    .CLK(dco_clk),
    .D(_02976_),
    .Q( execution_unit_0.inst_sext_5_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10205_ (
    .CLK(dco_clk),
    .D(_02977_),
    .Q( execution_unit_0.inst_sext_6_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10206_ (
    .CLK(dco_clk),
    .D(_02978_),
    .Q( execution_unit_0.inst_sext_7_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10207_ (
    .CLK(dco_clk),
    .D(_02979_),
    .Q( execution_unit_0.inst_sext_8_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10208_ (
    .CLK(dco_clk),
    .D(_02980_),
    .Q( execution_unit_0.inst_sext_9_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10209_ (
    .CLK(dco_clk),
    .D(_02981_),
    .Q( execution_unit_0.inst_sext_10_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10210_ (
    .CLK(dco_clk),
    .D(_02982_),
    .Q( execution_unit_0.inst_sext_11_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10211_ (
    .CLK(dco_clk),
    .D(_02983_),
    .Q( execution_unit_0.inst_sext_12_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10212_ (
    .CLK(dco_clk),
    .D(_02984_),
    .Q( execution_unit_0.inst_sext_13_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10213_ (
    .CLK(dco_clk),
    .D(_02985_),
    .Q( execution_unit_0.inst_sext_14_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10214_ (
    .CLK(dco_clk),
    .D(_02986_),
    .Q( execution_unit_0.inst_sext_15_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10215_ (
    .CLK(dco_clk),
    .D(_02987_),
    .Q( execution_unit_0.inst_ad_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10216_ (
    .CLK(dco_clk),
    .D(_02988_),
    .Q( execution_unit_0.UNUSED_inst_ad_idx ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10217_ (
    .CLK(dco_clk),
    .D(_02989_),
    .Q( execution_unit_0.UNUSED_inst_ad_symb ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10218_ (
    .CLK(dco_clk),
    .D(_02990_),
    .Q( execution_unit_0.inst_ad_6_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10219_ (
    .CLK(dco_clk),
    .D(_02906_),
    .Q( dbg_0.cpu_stat_full_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10220_ (
    .CLK(dco_clk),
    .D( frontend_0.i_state_nxt_0_ ),
    .Q( frontend_0.i_state_0_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10221_ (
    .CLK(dco_clk),
    .D( frontend_0.i_state_nxt_1_ ),
    .Q( frontend_0.i_state_1_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10222_ (
    .CLK(dco_clk),
    .D( frontend_0.i_state_nxt_2_ ),
    .Q( frontend_0.i_state_2_ ),
    .R(_02907_),
    .S(1'h1)
  );
  DFFSR _10223_ (
    .CLK(dco_clk),
    .D(_02991_),
    .Q( execution_unit_0.inst_irq_rst ),
    .R(1'h1),
    .S(_02907_)
  );
  DFFSR _10224_ (
    .CLK(dco_clk),
    .D(_02992_),
    .Q( frontend_0.irq_addr_1_ ),
    .R(1'h1),
    .S(_02907_)
  );
  DFFSR _10225_ (
    .CLK(dco_clk),
    .D(_02993_),
    .Q( frontend_0.irq_addr_2_ ),
    .R(1'h1),
    .S(_02907_)
  );
  DFFSR _10226_ (
    .CLK(dco_clk),
    .D(_02994_),
    .Q( frontend_0.irq_addr_3_ ),
    .R(1'h1),
    .S(_02907_)
  );
  DFFSR _10227_ (
    .CLK(dco_clk),
    .D(_02995_),
    .Q( frontend_0.irq_addr_4_ ),
    .R(1'h1),
    .S(_02907_)
  );
  INVX1 _10228_ (
    .A( dbg_0.cpu_stat_full_0_ ),
    .Y(_03737_)
  );
  INVX1 _10229_ (
    .A( dbg_0.UNUSED_eu_mb_wr_0_ ),
    .Y(_03738_)
  );
  INVX1 _10230_ (
    .A( dbg_0.dbg_mem_wr_0_ ),
    .Y(_03739_)
  );
  INVX1 _10231_ (
    .A( dbg_0.dbg_mem_addr_13_ ),
    .Y(_03740_)
  );
  INVX1 _10232_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .Y(_03741_)
  );
  INVX1 _10233_ (
    .A( dbg_0.dbg_mem_addr_10_ ),
    .Y(_03742_)
  );
  INVX1 _10234_ (
    .A( dbg_0.dbg_mem_addr_9_ ),
    .Y(_03743_)
  );
  INVX1 _10235_ (
    .A( dbg_0.dbg_mem_addr_12_ ),
    .Y(_03744_)
  );
  INVX1 _10236_ (
    .A( dbg_0.dbg_mem_addr_11_ ),
    .Y(_03745_)
  );
  INVX1 _10237_ (
    .A( dbg_0.dbg_mem_addr_2_ ),
    .Y(_03746_)
  );
  INVX1 _10238_ (
    .A( dbg_0.dbg_mem_addr_1_ ),
    .Y(_03747_)
  );
  INVX1 _10239_ (
    .A( dbg_0.dbg_mem_addr_4_ ),
    .Y(_03748_)
  );
  INVX1 _10240_ (
    .A( dbg_0.dbg_mem_addr_3_ ),
    .Y(_03749_)
  );
  INVX1 _10241_ (
    .A( dbg_0.dbg_mem_addr_6_ ),
    .Y(_03750_)
  );
  INVX1 _10242_ (
    .A( dbg_0.dbg_mem_addr_5_ ),
    .Y(_03751_)
  );
  INVX1 _10243_ (
    .A( dbg_0.dbg_mem_addr_8_ ),
    .Y(_03752_)
  );
  INVX1 _10244_ (
    .A( dbg_0.dbg_mem_addr_7_ ),
    .Y(_03753_)
  );
  INVX1 _10245_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .Y(_03754_)
  );
  INVX1 _10246_ (
    .A( dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_03755_)
  );
  INVX1 _10247_ (
    .A( dbg_0.UNUSED_eu_mab_10_ ),
    .Y(_03756_)
  );
  INVX1 _10248_ (
    .A( dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_03757_)
  );
  INVX1 _10249_ (
    .A( dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_03758_)
  );
  INVX1 _10250_ (
    .A( dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_03759_)
  );
  INVX1 _10251_ (
    .A( dbg_0.UNUSED_eu_mab_6_ ),
    .Y(_03760_)
  );
  INVX1 _10252_ (
    .A( dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_03761_)
  );
  INVX1 _10253_ (
    .A( dbg_0.UNUSED_eu_mab_8_ ),
    .Y(_03762_)
  );
  INVX1 _10254_ (
    .A( dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_03763_)
  );
  INVX1 _10255_ (
    .A( dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_03764_)
  );
  INVX1 _10256_ (
    .A( dbg_0.UNUSED_eu_mab_1_ ),
    .Y(_03765_)
  );
  INVX1 _10257_ (
    .A( dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_03766_)
  );
  INVX1 _10258_ (
    .A( dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_03767_)
  );
  INVX1 _10259_ (
    .A( dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_03768_)
  );
  INVX1 _10260_ (
    .A( dbg_0.dbg_mem_wr_1_ ),
    .Y(_03769_)
  );
  INVX1 _10261_ (
    .A(_05677_),
    .Y(_03770_)
  );
  INVX1 _10262_ (
    .A( execution_unit_0.mdb_out_0_ ),
    .Y(_03771_)
  );
  INVX1 _10263_ (
    .A(_05684_),
    .Y(_03772_)
  );
  INVX1 _10264_ (
    .A( execution_unit_0.mdb_out_1_ ),
    .Y(_03773_)
  );
  INVX1 _10265_ (
    .A(_05685_),
    .Y(_03774_)
  );
  INVX1 _10266_ (
    .A( execution_unit_0.mdb_out_2_ ),
    .Y(_03775_)
  );
  INVX1 _10267_ (
    .A(_05686_),
    .Y(_03776_)
  );
  INVX1 _10268_ (
    .A( execution_unit_0.mdb_out_3_ ),
    .Y(_03777_)
  );
  INVX1 _10269_ (
    .A(_05687_),
    .Y(_03778_)
  );
  INVX1 _10270_ (
    .A( execution_unit_0.mdb_out_4_ ),
    .Y(_03779_)
  );
  INVX1 _10271_ (
    .A(_05688_),
    .Y(_03780_)
  );
  INVX1 _10272_ (
    .A( execution_unit_0.mdb_out_5_ ),
    .Y(_03781_)
  );
  INVX1 _10273_ (
    .A(_05689_),
    .Y(_03782_)
  );
  INVX1 _10274_ (
    .A( execution_unit_0.mdb_out_6_ ),
    .Y(_03783_)
  );
  INVX1 _10275_ (
    .A(_05690_),
    .Y(_03784_)
  );
  INVX1 _10276_ (
    .A( execution_unit_0.mdb_out_7_ ),
    .Y(_03785_)
  );
  INVX1 _10277_ (
    .A(_05691_),
    .Y(_03786_)
  );
  INVX1 _10278_ (
    .A( execution_unit_0.mdb_out_8_ ),
    .Y(_03787_)
  );
  INVX1 _10279_ (
    .A(_05692_),
    .Y(_03788_)
  );
  INVX1 _10280_ (
    .A( execution_unit_0.mdb_out_9_ ),
    .Y(_03789_)
  );
  INVX1 _10281_ (
    .A(_05678_),
    .Y(_03790_)
  );
  INVX1 _10282_ (
    .A( execution_unit_0.mdb_out_10_ ),
    .Y(_03791_)
  );
  INVX1 _10283_ (
    .A(_05679_),
    .Y(_03792_)
  );
  INVX1 _10284_ (
    .A( execution_unit_0.mdb_out_11_ ),
    .Y(_03793_)
  );
  INVX1 _10285_ (
    .A(_05680_),
    .Y(_03794_)
  );
  INVX1 _10286_ (
    .A( execution_unit_0.mdb_out_12_ ),
    .Y(_03795_)
  );
  INVX1 _10287_ (
    .A(_05681_),
    .Y(_03796_)
  );
  INVX1 _10288_ (
    .A( execution_unit_0.mdb_out_13_ ),
    .Y(_03797_)
  );
  INVX1 _10289_ (
    .A(_05682_),
    .Y(_03798_)
  );
  INVX1 _10290_ (
    .A( execution_unit_0.mdb_out_14_ ),
    .Y(_03799_)
  );
  INVX1 _10291_ (
    .A(_05683_),
    .Y(_03800_)
  );
  INVX1 _10292_ (
    .A( execution_unit_0.mdb_out_15_ ),
    .Y(_03801_)
  );
  INVX1 _10293_ (
    .A(pmem_dout_0_),
    .Y(_03802_)
  );
  INVX1 _10294_ (
    .A(pmem_dout_1_),
    .Y(_03803_)
  );
  INVX1 _10295_ (
    .A(pmem_dout_2_),
    .Y(_03804_)
  );
  INVX1 _10296_ (
    .A(pmem_dout_3_),
    .Y(_03805_)
  );
  INVX1 _10297_ (
    .A(pmem_dout_4_),
    .Y(_03806_)
  );
  INVX1 _10298_ (
    .A(pmem_dout_5_),
    .Y(_03807_)
  );
  INVX1 _10299_ (
    .A(pmem_dout_6_),
    .Y(_03808_)
  );
  INVX1 _10300_ (
    .A(pmem_dout_7_),
    .Y(_03809_)
  );
  INVX1 _10301_ (
    .A(pmem_dout_8_),
    .Y(_03810_)
  );
  INVX1 _10302_ (
    .A(pmem_dout_9_),
    .Y(_03811_)
  );
  INVX1 _10303_ (
    .A(pmem_dout_10_),
    .Y(_03812_)
  );
  INVX1 _10304_ (
    .A(pmem_dout_11_),
    .Y(_03813_)
  );
  INVX1 _10305_ (
    .A(pmem_dout_12_),
    .Y(_03814_)
  );
  INVX1 _10306_ (
    .A(pmem_dout_13_),
    .Y(_03815_)
  );
  INVX1 _10307_ (
    .A(pmem_dout_14_),
    .Y(_03816_)
  );
  INVX1 _10308_ (
    .A(pmem_dout_15_),
    .Y(_03817_)
  );
  INVX1 _10309_ (
    .A(_05695_),
    .Y(_03719_)
  );
  NAND2X1 _10310_ (
    .A( frontend_0.mb_en ),
    .B( execution_unit_0.pc_nxt_15_ ),
    .Y(_03818_)
  );
  INVX1 _10311_ (
    .A(_03818_),
    .Y( mem_backbone_0.fe_pmem_en )
  );
  NAND2X1 _10312_ (
    .A( dbg_0.UNUSED_eu_mab_14_ ),
    .B( dbg_0.UNUSED_eu_mb_en ),
    .Y(_03819_)
  );
  NOR2X1 _10313_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B(_03819_),
    .Y(_03820_)
  );
  NAND3X1 _10314_ (
    .A( dbg_0.dbg_mem_addr_14_ ),
    .B(_03754_),
    .C( dbg_0.dbg_mem_en ),
    .Y(_03821_)
  );
  NOR2X1 _10315_ (
    .A(_03820_),
    .B(_03821_),
    .Y(_03822_)
  );
  MUX2X1 _10316_ (
    .A( dbg_0.dbg_mem_wr_0_ ),
    .B( dbg_0.UNUSED_eu_mb_wr_0_ ),
    .S(_03822_),
    .Y(_05614_)
  );
  MUX2X1 _10317_ (
    .A( dbg_0.dbg_mem_wr_1_ ),
    .B( dbg_0.UNUSED_eu_mb_wr_1_ ),
    .S(_03822_),
    .Y(_05615_)
  );
  MUX2X1 _10318_ (
    .A(_03747_),
    .B(_03765_),
    .S(_03822_),
    .Y(_05584_)
  );
  MUX2X1 _10319_ (
    .A(_03746_),
    .B(_03764_),
    .S(_03822_),
    .Y(_05588_)
  );
  MUX2X1 _10320_ (
    .A(_03749_),
    .B(_03767_),
    .S(_03822_),
    .Y(_05589_)
  );
  MUX2X1 _10321_ (
    .A(_03748_),
    .B(_03766_),
    .S(_03822_),
    .Y(_05590_)
  );
  MUX2X1 _10322_ (
    .A(_03751_),
    .B(_03761_),
    .S(_03822_),
    .Y(_05591_)
  );
  MUX2X1 _10323_ (
    .A(_03750_),
    .B(_03760_),
    .S(_03822_),
    .Y(_05592_)
  );
  MUX2X1 _10324_ (
    .A(_03753_),
    .B(_03763_),
    .S(_03822_),
    .Y(_05593_)
  );
  MUX2X1 _10325_ (
    .A(_03752_),
    .B(_03762_),
    .S(_03822_),
    .Y(_05594_)
  );
  MUX2X1 _10326_ (
    .A(_03743_),
    .B(_03757_),
    .S(_03822_),
    .Y(_05595_)
  );
  MUX2X1 _10327_ (
    .A(_03742_),
    .B(_03756_),
    .S(_03822_),
    .Y(_05596_)
  );
  MUX2X1 _10328_ (
    .A(_03745_),
    .B(_03759_),
    .S(_03822_),
    .Y(_05585_)
  );
  MUX2X1 _10329_ (
    .A(_03744_),
    .B(_03758_),
    .S(_03822_),
    .Y(_05586_)
  );
  MUX2X1 _10330_ (
    .A(_03740_),
    .B(_03755_),
    .S(_03822_),
    .Y(_05587_)
  );
  MUX2X1 _10331_ (
    .A(_03770_),
    .B(_03771_),
    .S(_03822_),
    .Y(_05598_)
  );
  MUX2X1 _10332_ (
    .A(_03772_),
    .B(_03773_),
    .S(_03822_),
    .Y(_05605_)
  );
  MUX2X1 _10333_ (
    .A(_03774_),
    .B(_03775_),
    .S(_03822_),
    .Y(_05606_)
  );
  MUX2X1 _10334_ (
    .A(_03776_),
    .B(_03777_),
    .S(_03822_),
    .Y(_05607_)
  );
  MUX2X1 _10335_ (
    .A(_03778_),
    .B(_03779_),
    .S(_03822_),
    .Y(_05608_)
  );
  MUX2X1 _10336_ (
    .A(_03780_),
    .B(_03781_),
    .S(_03822_),
    .Y(_05609_)
  );
  MUX2X1 _10337_ (
    .A(_03782_),
    .B(_03783_),
    .S(_03822_),
    .Y(_05610_)
  );
  MUX2X1 _10338_ (
    .A(_03784_),
    .B(_03785_),
    .S(_03822_),
    .Y(_05611_)
  );
  MUX2X1 _10339_ (
    .A(_03786_),
    .B(_03787_),
    .S(_03822_),
    .Y(_05612_)
  );
  MUX2X1 _10340_ (
    .A(_03788_),
    .B(_03789_),
    .S(_03822_),
    .Y(_05613_)
  );
  MUX2X1 _10341_ (
    .A(_03790_),
    .B(_03791_),
    .S(_03822_),
    .Y(_05599_)
  );
  MUX2X1 _10342_ (
    .A(_03792_),
    .B(_03793_),
    .S(_03822_),
    .Y(_05600_)
  );
  MUX2X1 _10343_ (
    .A(_03794_),
    .B(_03795_),
    .S(_03822_),
    .Y(_05601_)
  );
  MUX2X1 _10344_ (
    .A(_03796_),
    .B(_03797_),
    .S(_03822_),
    .Y(_05602_)
  );
  MUX2X1 _10345_ (
    .A(_03798_),
    .B(_03799_),
    .S(_03822_),
    .Y(_05603_)
  );
  MUX2X1 _10346_ (
    .A(_03800_),
    .B(_03801_),
    .S(_03822_),
    .Y(_05604_)
  );
  OR2X1 _10347_ (
    .A( dbg_0.UNUSED_eu_mb_wr_0_ ),
    .B( dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_03823_)
  );
  NAND2X1 _10348_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B( dbg_0.UNUSED_eu_mb_en ),
    .Y(_03824_)
  );
  NOR2X1 _10349_ (
    .A(_03823_),
    .B(_03824_),
    .Y( mem_backbone_0.eu_pmem_en )
  );
  OAI21X1 _10350_ (
    .A(_03823_),
    .B(_03824_),
    .C(_03818_),
    .Y(_03825_)
  );
  NAND2X1 _10351_ (
    .A( dbg_0.dbg_mem_addr_15_ ),
    .B( dbg_0.dbg_mem_en ),
    .Y(_03826_)
  );
  NOR2X1 _10352_ (
    .A(_03825_),
    .B(_03826_),
    .Y( mem_backbone_0.ext_pmem_en )
  );
  NAND2X1 _10353_ (
    .A( dbg_0.dbg_mem_wr_0_ ),
    .B( mem_backbone_0.ext_pmem_en ),
    .Y(_05693_)
  );
  NAND2X1 _10354_ (
    .A( dbg_0.dbg_mem_wr_1_ ),
    .B( mem_backbone_0.ext_pmem_en ),
    .Y(_05694_)
  );
  MUX2X1 _10355_ (
    .A( dbg_0.UNUSED_eu_mab_1_ ),
    .B( execution_unit_0.pc_nxt_1_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03827_)
  );
  MUX2X1 _10356_ (
    .A(_03747_),
    .B(_03827_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05662_)
  );
  MUX2X1 _10357_ (
    .A( dbg_0.UNUSED_eu_mab_2_ ),
    .B( execution_unit_0.pc_nxt_2_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03828_)
  );
  MUX2X1 _10358_ (
    .A(_03746_),
    .B(_03828_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05667_)
  );
  MUX2X1 _10359_ (
    .A( dbg_0.UNUSED_eu_mab_3_ ),
    .B( execution_unit_0.pc_nxt_3_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03829_)
  );
  MUX2X1 _10360_ (
    .A(_03749_),
    .B(_03829_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05668_)
  );
  MUX2X1 _10361_ (
    .A( dbg_0.UNUSED_eu_mab_4_ ),
    .B( execution_unit_0.pc_nxt_4_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03830_)
  );
  MUX2X1 _10362_ (
    .A(_03748_),
    .B(_03830_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05669_)
  );
  MUX2X1 _10363_ (
    .A( dbg_0.UNUSED_eu_mab_5_ ),
    .B( execution_unit_0.pc_nxt_5_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03831_)
  );
  MUX2X1 _10364_ (
    .A(_03751_),
    .B(_03831_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05670_)
  );
  MUX2X1 _10365_ (
    .A( dbg_0.UNUSED_eu_mab_6_ ),
    .B( execution_unit_0.pc_nxt_6_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03832_)
  );
  MUX2X1 _10366_ (
    .A(_03750_),
    .B(_03832_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05671_)
  );
  MUX2X1 _10367_ (
    .A( dbg_0.UNUSED_eu_mab_7_ ),
    .B( execution_unit_0.pc_nxt_7_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03833_)
  );
  MUX2X1 _10368_ (
    .A(_03753_),
    .B(_03833_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05672_)
  );
  MUX2X1 _10369_ (
    .A( dbg_0.UNUSED_eu_mab_8_ ),
    .B( execution_unit_0.pc_nxt_8_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03834_)
  );
  MUX2X1 _10370_ (
    .A(_03752_),
    .B(_03834_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05673_)
  );
  MUX2X1 _10371_ (
    .A( dbg_0.UNUSED_eu_mab_9_ ),
    .B( execution_unit_0.pc_nxt_9_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03835_)
  );
  MUX2X1 _10372_ (
    .A(_03743_),
    .B(_03835_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05674_)
  );
  MUX2X1 _10373_ (
    .A( dbg_0.UNUSED_eu_mab_10_ ),
    .B( execution_unit_0.pc_nxt_10_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03836_)
  );
  MUX2X1 _10374_ (
    .A(_03742_),
    .B(_03836_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05675_)
  );
  MUX2X1 _10375_ (
    .A( dbg_0.UNUSED_eu_mab_11_ ),
    .B( execution_unit_0.pc_nxt_11_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03837_)
  );
  MUX2X1 _10376_ (
    .A(_03745_),
    .B(_03837_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05663_)
  );
  MUX2X1 _10377_ (
    .A( dbg_0.UNUSED_eu_mab_12_ ),
    .B( execution_unit_0.pc_nxt_12_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03838_)
  );
  MUX2X1 _10378_ (
    .A(_03744_),
    .B(_03838_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05664_)
  );
  MUX2X1 _10379_ (
    .A( dbg_0.UNUSED_eu_mab_13_ ),
    .B( execution_unit_0.pc_nxt_13_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03839_)
  );
  MUX2X1 _10380_ (
    .A(_03740_),
    .B(_03839_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05665_)
  );
  MUX2X1 _10381_ (
    .A( dbg_0.UNUSED_eu_mab_14_ ),
    .B( execution_unit_0.pc_nxt_14_ ),
    .S( mem_backbone_0.eu_pmem_en ),
    .Y(_03840_)
  );
  MUX2X1 _10382_ (
    .A(_03741_),
    .B(_03840_),
    .S( mem_backbone_0.ext_pmem_en ),
    .Y(_05666_)
  );
  NOR2X1 _10383_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B( dbg_0.UNUSED_eu_mab_14_ ),
    .Y(_03841_)
  );
  NAND2X1 _10384_ (
    .A( dbg_0.UNUSED_eu_mb_en ),
    .B(_03841_),
    .Y(_03842_)
  );
  INVX1 _10385_ (
    .A(_03842_),
    .Y( mem_backbone_0.eu_per_en )
  );
  NAND3X1 _10386_ (
    .A(_03741_),
    .B(_03754_),
    .C( dbg_0.dbg_mem_en ),
    .Y(_03843_)
  );
  NOR2X1 _10387_ (
    .A( mem_backbone_0.eu_per_en ),
    .B(_03843_),
    .Y( mem_backbone_0.ext_per_en )
  );
  MUX2X1 _10388_ (
    .A(_03739_),
    .B(_03738_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05660_)
  );
  MUX2X1 _10389_ (
    .A(_03769_),
    .B(_03768_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05661_)
  );
  MUX2X1 _10390_ (
    .A(_03747_),
    .B(_03765_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05630_)
  );
  MUX2X1 _10391_ (
    .A(_03746_),
    .B(_03764_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05634_)
  );
  MUX2X1 _10392_ (
    .A(_03749_),
    .B(_03767_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05635_)
  );
  MUX2X1 _10393_ (
    .A(_03748_),
    .B(_03766_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05636_)
  );
  MUX2X1 _10394_ (
    .A(_03751_),
    .B(_03761_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05637_)
  );
  MUX2X1 _10395_ (
    .A(_03750_),
    .B(_03760_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05638_)
  );
  MUX2X1 _10396_ (
    .A(_03753_),
    .B(_03763_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05639_)
  );
  MUX2X1 _10397_ (
    .A(_03752_),
    .B(_03762_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05640_)
  );
  MUX2X1 _10398_ (
    .A(_03743_),
    .B(_03757_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05641_)
  );
  MUX2X1 _10399_ (
    .A(_03742_),
    .B(_03756_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05642_)
  );
  MUX2X1 _10400_ (
    .A(_03745_),
    .B(_03759_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05631_)
  );
  MUX2X1 _10401_ (
    .A(_03744_),
    .B(_03758_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05632_)
  );
  MUX2X1 _10402_ (
    .A(_03740_),
    .B(_03755_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05633_)
  );
  MUX2X1 _10403_ (
    .A(_03770_),
    .B(_03771_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05643_)
  );
  MUX2X1 _10404_ (
    .A(_03772_),
    .B(_03773_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05650_)
  );
  MUX2X1 _10405_ (
    .A(_03774_),
    .B(_03775_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05651_)
  );
  MUX2X1 _10406_ (
    .A(_03776_),
    .B(_03777_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05652_)
  );
  MUX2X1 _10407_ (
    .A(_03778_),
    .B(_03779_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05653_)
  );
  MUX2X1 _10408_ (
    .A(_03780_),
    .B(_03781_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05654_)
  );
  MUX2X1 _10409_ (
    .A(_03782_),
    .B(_03783_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05655_)
  );
  MUX2X1 _10410_ (
    .A(_03784_),
    .B(_03785_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05656_)
  );
  MUX2X1 _10411_ (
    .A(_03786_),
    .B(_03787_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05657_)
  );
  MUX2X1 _10412_ (
    .A(_03788_),
    .B(_03789_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05658_)
  );
  MUX2X1 _10413_ (
    .A(_03790_),
    .B(_03791_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05644_)
  );
  MUX2X1 _10414_ (
    .A(_03792_),
    .B(_03793_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05645_)
  );
  MUX2X1 _10415_ (
    .A(_03794_),
    .B(_03795_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05646_)
  );
  MUX2X1 _10416_ (
    .A(_03796_),
    .B(_03797_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05647_)
  );
  MUX2X1 _10417_ (
    .A(_03798_),
    .B(_03799_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05648_)
  );
  MUX2X1 _10418_ (
    .A(_03800_),
    .B(_03801_),
    .S( mem_backbone_0.ext_per_en ),
    .Y(_05649_)
  );
  NAND2X1 _10419_ (
    .A( mem_backbone_0.pmem_dout_bckup_0_ ),
    .B( mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_03844_)
  );
  OAI21X1 _10420_ (
    .A(_03802_),
    .B( mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_03844_),
    .Y( dbg_0.fe_mdb_in_0_ )
  );
  NAND2X1 _10421_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_1_ ),
    .Y(_03845_)
  );
  OAI21X1 _10422_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03803_),
    .C(_03845_),
    .Y( dbg_0.fe_mdb_in_1_ )
  );
  NAND2X1 _10423_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_2_ ),
    .Y(_03846_)
  );
  OAI21X1 _10424_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03804_),
    .C(_03846_),
    .Y( dbg_0.fe_mdb_in_2_ )
  );
  NAND2X1 _10425_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_3_ ),
    .Y(_03847_)
  );
  OAI21X1 _10426_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03805_),
    .C(_03847_),
    .Y( dbg_0.fe_mdb_in_3_ )
  );
  NAND2X1 _10427_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_4_ ),
    .Y(_03848_)
  );
  OAI21X1 _10428_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03806_),
    .C(_03848_),
    .Y( dbg_0.fe_mdb_in_4_ )
  );
  NAND2X1 _10429_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_5_ ),
    .Y(_03849_)
  );
  OAI21X1 _10430_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03807_),
    .C(_03849_),
    .Y( dbg_0.fe_mdb_in_5_ )
  );
  NAND2X1 _10431_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_6_ ),
    .Y(_03850_)
  );
  OAI21X1 _10432_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03808_),
    .C(_03850_),
    .Y( dbg_0.fe_mdb_in_6_ )
  );
  NAND2X1 _10433_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_7_ ),
    .Y(_03851_)
  );
  OAI21X1 _10434_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03809_),
    .C(_03851_),
    .Y( dbg_0.fe_mdb_in_7_ )
  );
  NAND2X1 _10435_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_8_ ),
    .Y(_03852_)
  );
  OAI21X1 _10436_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03810_),
    .C(_03852_),
    .Y( dbg_0.fe_mdb_in_8_ )
  );
  NAND2X1 _10437_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_9_ ),
    .Y(_03853_)
  );
  OAI21X1 _10438_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03811_),
    .C(_03853_),
    .Y( dbg_0.fe_mdb_in_9_ )
  );
  NAND2X1 _10439_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_10_ ),
    .Y(_03854_)
  );
  OAI21X1 _10440_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03812_),
    .C(_03854_),
    .Y( dbg_0.fe_mdb_in_10_ )
  );
  NAND2X1 _10441_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_11_ ),
    .Y(_03855_)
  );
  OAI21X1 _10442_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03813_),
    .C(_03855_),
    .Y( dbg_0.fe_mdb_in_11_ )
  );
  NAND2X1 _10443_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_12_ ),
    .Y(_03856_)
  );
  OAI21X1 _10444_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03814_),
    .C(_03856_),
    .Y( dbg_0.fe_mdb_in_12_ )
  );
  NAND2X1 _10445_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_13_ ),
    .Y(_03857_)
  );
  OAI21X1 _10446_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03815_),
    .C(_03857_),
    .Y( dbg_0.fe_mdb_in_13_ )
  );
  NAND2X1 _10447_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_14_ ),
    .Y(_03858_)
  );
  OAI21X1 _10448_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03816_),
    .C(_03858_),
    .Y( dbg_0.fe_mdb_in_14_ )
  );
  NAND2X1 _10449_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B( mem_backbone_0.pmem_dout_bckup_15_ ),
    .Y(_03859_)
  );
  OAI21X1 _10450_ (
    .A( mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_03817_),
    .C(_03859_),
    .Y( dbg_0.fe_mdb_in_15_ )
  );
  MUX2X1 _10451_ (
    .A( mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03860_)
  );
  NAND2X1 _10452_ (
    .A(pmem_dout_0_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03861_)
  );
  OAI21X1 _10453_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03860_),
    .C(_03861_),
    .Y( execution_unit_0.mdb_in_0_ )
  );
  MUX2X1 _10454_ (
    .A( mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03862_)
  );
  NAND2X1 _10455_ (
    .A(pmem_dout_1_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03863_)
  );
  OAI21X1 _10456_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03862_),
    .C(_03863_),
    .Y( execution_unit_0.mdb_in_1_ )
  );
  MUX2X1 _10457_ (
    .A( mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03864_)
  );
  NAND2X1 _10458_ (
    .A(pmem_dout_2_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03865_)
  );
  OAI21X1 _10459_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03864_),
    .C(_03865_),
    .Y( execution_unit_0.mdb_in_2_ )
  );
  MUX2X1 _10460_ (
    .A( mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03866_)
  );
  NAND2X1 _10461_ (
    .A(pmem_dout_3_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03867_)
  );
  OAI21X1 _10462_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03866_),
    .C(_03867_),
    .Y( execution_unit_0.mdb_in_3_ )
  );
  MUX2X1 _10463_ (
    .A( mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03868_)
  );
  NAND2X1 _10464_ (
    .A(pmem_dout_4_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03869_)
  );
  OAI21X1 _10465_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03868_),
    .C(_03869_),
    .Y( execution_unit_0.mdb_in_4_ )
  );
  MUX2X1 _10466_ (
    .A( mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03870_)
  );
  NAND2X1 _10467_ (
    .A(pmem_dout_5_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03871_)
  );
  OAI21X1 _10468_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03870_),
    .C(_03871_),
    .Y( execution_unit_0.mdb_in_5_ )
  );
  MUX2X1 _10469_ (
    .A( mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03872_)
  );
  NAND2X1 _10470_ (
    .A(pmem_dout_6_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03873_)
  );
  OAI21X1 _10471_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03872_),
    .C(_03873_),
    .Y( execution_unit_0.mdb_in_6_ )
  );
  MUX2X1 _10472_ (
    .A( mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03874_)
  );
  NAND2X1 _10473_ (
    .A(pmem_dout_7_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03875_)
  );
  OAI21X1 _10474_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03874_),
    .C(_03875_),
    .Y( execution_unit_0.mdb_in_7_ )
  );
  MUX2X1 _10475_ (
    .A( mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03876_)
  );
  NAND2X1 _10476_ (
    .A(pmem_dout_8_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03877_)
  );
  OAI21X1 _10477_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03876_),
    .C(_03877_),
    .Y( execution_unit_0.mdb_in_8_ )
  );
  MUX2X1 _10478_ (
    .A( mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03878_)
  );
  NAND2X1 _10479_ (
    .A(pmem_dout_9_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03879_)
  );
  OAI21X1 _10480_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03878_),
    .C(_03879_),
    .Y( execution_unit_0.mdb_in_9_ )
  );
  MUX2X1 _10481_ (
    .A( mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03880_)
  );
  NAND2X1 _10482_ (
    .A(pmem_dout_10_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03881_)
  );
  OAI21X1 _10483_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03880_),
    .C(_03881_),
    .Y( execution_unit_0.mdb_in_10_ )
  );
  MUX2X1 _10484_ (
    .A( mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03882_)
  );
  NAND2X1 _10485_ (
    .A(pmem_dout_11_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03883_)
  );
  OAI21X1 _10486_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03882_),
    .C(_03883_),
    .Y( execution_unit_0.mdb_in_11_ )
  );
  MUX2X1 _10487_ (
    .A( mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03884_)
  );
  NAND2X1 _10488_ (
    .A(pmem_dout_12_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03885_)
  );
  OAI21X1 _10489_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03884_),
    .C(_03885_),
    .Y( execution_unit_0.mdb_in_12_ )
  );
  MUX2X1 _10490_ (
    .A( mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03886_)
  );
  NAND2X1 _10491_ (
    .A(pmem_dout_13_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03887_)
  );
  OAI21X1 _10492_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03886_),
    .C(_03887_),
    .Y( execution_unit_0.mdb_in_13_ )
  );
  MUX2X1 _10493_ (
    .A( mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03888_)
  );
  NAND2X1 _10494_ (
    .A(pmem_dout_14_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03889_)
  );
  OAI21X1 _10495_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03888_),
    .C(_03889_),
    .Y( execution_unit_0.mdb_in_14_ )
  );
  MUX2X1 _10496_ (
    .A( mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_03890_)
  );
  NAND2X1 _10497_ (
    .A(pmem_dout_15_),
    .B( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_03891_)
  );
  OAI21X1 _10498_ (
    .A( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_03890_),
    .C(_03891_),
    .Y( execution_unit_0.mdb_in_15_ )
  );
  MUX2X1 _10499_ (
    .A( mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03892_)
  );
  NAND2X1 _10500_ (
    .A(pmem_dout_0_),
    .B(_03718_),
    .Y(_03893_)
  );
  OAI21X1 _10501_ (
    .A(_03718_),
    .B(_03892_),
    .C(_03893_),
    .Y( dbg_0.dbg_mem_din_0_ )
  );
  MUX2X1 _10502_ (
    .A( mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03894_)
  );
  NAND2X1 _10503_ (
    .A(pmem_dout_1_),
    .B(_03718_),
    .Y(_03895_)
  );
  OAI21X1 _10504_ (
    .A(_03718_),
    .B(_03894_),
    .C(_03895_),
    .Y( dbg_0.dbg_mem_din_1_ )
  );
  MUX2X1 _10505_ (
    .A( mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03896_)
  );
  NAND2X1 _10506_ (
    .A(pmem_dout_2_),
    .B(_03718_),
    .Y(_03897_)
  );
  OAI21X1 _10507_ (
    .A(_03718_),
    .B(_03896_),
    .C(_03897_),
    .Y( dbg_0.dbg_mem_din_2_ )
  );
  MUX2X1 _10508_ (
    .A( mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03898_)
  );
  NAND2X1 _10509_ (
    .A(pmem_dout_3_),
    .B(_03718_),
    .Y(_03899_)
  );
  OAI21X1 _10510_ (
    .A(_03718_),
    .B(_03898_),
    .C(_03899_),
    .Y( dbg_0.dbg_mem_din_3_ )
  );
  MUX2X1 _10511_ (
    .A( mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03900_)
  );
  NAND2X1 _10512_ (
    .A(pmem_dout_4_),
    .B(_03718_),
    .Y(_03901_)
  );
  OAI21X1 _10513_ (
    .A(_03718_),
    .B(_03900_),
    .C(_03901_),
    .Y( dbg_0.dbg_mem_din_4_ )
  );
  MUX2X1 _10514_ (
    .A( mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03902_)
  );
  NAND2X1 _10515_ (
    .A(pmem_dout_5_),
    .B(_03718_),
    .Y(_03903_)
  );
  OAI21X1 _10516_ (
    .A(_03718_),
    .B(_03902_),
    .C(_03903_),
    .Y( dbg_0.dbg_mem_din_5_ )
  );
  MUX2X1 _10517_ (
    .A( mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03904_)
  );
  NAND2X1 _10518_ (
    .A(pmem_dout_6_),
    .B(_03718_),
    .Y(_03905_)
  );
  OAI21X1 _10519_ (
    .A(_03718_),
    .B(_03904_),
    .C(_03905_),
    .Y( dbg_0.dbg_mem_din_6_ )
  );
  MUX2X1 _10520_ (
    .A( mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03906_)
  );
  NAND2X1 _10521_ (
    .A(pmem_dout_7_),
    .B(_03718_),
    .Y(_03907_)
  );
  OAI21X1 _10522_ (
    .A(_03718_),
    .B(_03906_),
    .C(_03907_),
    .Y( dbg_0.dbg_mem_din_7_ )
  );
  MUX2X1 _10523_ (
    .A( mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03908_)
  );
  NAND2X1 _10524_ (
    .A(pmem_dout_8_),
    .B(_03718_),
    .Y(_03909_)
  );
  OAI21X1 _10525_ (
    .A(_03718_),
    .B(_03908_),
    .C(_03909_),
    .Y( dbg_0.dbg_mem_din_8_ )
  );
  MUX2X1 _10526_ (
    .A( mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03910_)
  );
  NAND2X1 _10527_ (
    .A(pmem_dout_9_),
    .B(_03718_),
    .Y(_03911_)
  );
  OAI21X1 _10528_ (
    .A(_03718_),
    .B(_03910_),
    .C(_03911_),
    .Y( dbg_0.dbg_mem_din_9_ )
  );
  MUX2X1 _10529_ (
    .A( mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03912_)
  );
  NAND2X1 _10530_ (
    .A(pmem_dout_10_),
    .B(_03718_),
    .Y(_03913_)
  );
  OAI21X1 _10531_ (
    .A(_03718_),
    .B(_03912_),
    .C(_03913_),
    .Y( dbg_0.dbg_mem_din_10_ )
  );
  MUX2X1 _10532_ (
    .A( mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03914_)
  );
  NAND2X1 _10533_ (
    .A(pmem_dout_11_),
    .B(_03718_),
    .Y(_03915_)
  );
  OAI21X1 _10534_ (
    .A(_03718_),
    .B(_03914_),
    .C(_03915_),
    .Y( dbg_0.dbg_mem_din_11_ )
  );
  MUX2X1 _10535_ (
    .A( mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03916_)
  );
  NAND2X1 _10536_ (
    .A(pmem_dout_12_),
    .B(_03718_),
    .Y(_03917_)
  );
  OAI21X1 _10537_ (
    .A(_03718_),
    .B(_03916_),
    .C(_03917_),
    .Y( dbg_0.dbg_mem_din_12_ )
  );
  MUX2X1 _10538_ (
    .A( mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03918_)
  );
  NAND2X1 _10539_ (
    .A(pmem_dout_13_),
    .B(_03718_),
    .Y(_03919_)
  );
  OAI21X1 _10540_ (
    .A(_03718_),
    .B(_03918_),
    .C(_03919_),
    .Y( dbg_0.dbg_mem_din_13_ )
  );
  MUX2X1 _10541_ (
    .A( mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03920_)
  );
  NAND2X1 _10542_ (
    .A(pmem_dout_14_),
    .B(_03718_),
    .Y(_03921_)
  );
  OAI21X1 _10543_ (
    .A(_03718_),
    .B(_03920_),
    .C(_03921_),
    .Y( dbg_0.dbg_mem_din_14_ )
  );
  MUX2X1 _10544_ (
    .A( mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S( mem_backbone_0.ext_mem_din_sel ),
    .Y(_03922_)
  );
  NAND2X1 _10545_ (
    .A(pmem_dout_15_),
    .B(_03718_),
    .Y(_03923_)
  );
  OAI21X1 _10546_ (
    .A(_03718_),
    .B(_03922_),
    .C(_03923_),
    .Y( dbg_0.dbg_mem_din_15_ )
  );
  OAI21X1 _10547_ (
    .A( dbg_0.UNUSED_eu_mab_15_ ),
    .B(_03819_),
    .C(_03821_),
    .Y(_03924_)
  );
  INVX1 _10548_ (
    .A(_03924_),
    .Y(_05597_)
  );
  NOR2X1 _10549_ (
    .A(_03825_),
    .B( mem_backbone_0.ext_pmem_en ),
    .Y(_05676_)
  );
  AND2X1 _10550_ (
    .A( mem_backbone_0.fe_pmem_en ),
    .B( mem_backbone_0.eu_pmem_en ),
    .Y( frontend_0.fe_pmem_wait )
  );
  NAND2X1 _10551_ (
    .A(_03842_),
    .B(_03843_),
    .Y(_05659_)
  );
  NAND3X1 _10552_ (
    .A( mem_backbone_0.fe_pmem_en_dly ),
    .B(_03737_),
    .C(_03818_),
    .Y(_03925_)
  );
  MUX2X1 _10553_ (
    .A( mem_backbone_0.pmem_dout_bckup_0_ ),
    .B(pmem_dout_0_),
    .S(_03925_),
    .Y(_03926_)
  );
  INVX1 _10554_ (
    .A(_03926_),
    .Y(_03720_)
  );
  MUX2X1 _10555_ (
    .A( mem_backbone_0.pmem_dout_bckup_1_ ),
    .B(pmem_dout_1_),
    .S(_03925_),
    .Y(_03927_)
  );
  INVX1 _10556_ (
    .A(_03927_),
    .Y(_03721_)
  );
  MUX2X1 _10557_ (
    .A( mem_backbone_0.pmem_dout_bckup_2_ ),
    .B(pmem_dout_2_),
    .S(_03925_),
    .Y(_03928_)
  );
  INVX1 _10558_ (
    .A(_03928_),
    .Y(_03722_)
  );
  MUX2X1 _10559_ (
    .A( mem_backbone_0.pmem_dout_bckup_3_ ),
    .B(pmem_dout_3_),
    .S(_03925_),
    .Y(_03929_)
  );
  INVX1 _10560_ (
    .A(_03929_),
    .Y(_03723_)
  );
  MUX2X1 _10561_ (
    .A( mem_backbone_0.pmem_dout_bckup_4_ ),
    .B(pmem_dout_4_),
    .S(_03925_),
    .Y(_03930_)
  );
  INVX1 _10562_ (
    .A(_03930_),
    .Y(_03724_)
  );
  MUX2X1 _10563_ (
    .A( mem_backbone_0.pmem_dout_bckup_5_ ),
    .B(pmem_dout_5_),
    .S(_03925_),
    .Y(_03931_)
  );
  INVX1 _10564_ (
    .A(_03931_),
    .Y(_03725_)
  );
  MUX2X1 _10565_ (
    .A( mem_backbone_0.pmem_dout_bckup_6_ ),
    .B(pmem_dout_6_),
    .S(_03925_),
    .Y(_03932_)
  );
  INVX1 _10566_ (
    .A(_03932_),
    .Y(_03726_)
  );
  MUX2X1 _10567_ (
    .A( mem_backbone_0.pmem_dout_bckup_7_ ),
    .B(pmem_dout_7_),
    .S(_03925_),
    .Y(_03933_)
  );
  INVX1 _10568_ (
    .A(_03933_),
    .Y(_03727_)
  );
  MUX2X1 _10569_ (
    .A( mem_backbone_0.pmem_dout_bckup_8_ ),
    .B(pmem_dout_8_),
    .S(_03925_),
    .Y(_03934_)
  );
  INVX1 _10570_ (
    .A(_03934_),
    .Y(_03728_)
  );
  MUX2X1 _10571_ (
    .A( mem_backbone_0.pmem_dout_bckup_9_ ),
    .B(pmem_dout_9_),
    .S(_03925_),
    .Y(_03935_)
  );
  INVX1 _10572_ (
    .A(_03935_),
    .Y(_03729_)
  );
  MUX2X1 _10573_ (
    .A( mem_backbone_0.pmem_dout_bckup_10_ ),
    .B(pmem_dout_10_),
    .S(_03925_),
    .Y(_03936_)
  );
  INVX1 _10574_ (
    .A(_03936_),
    .Y(_03730_)
  );
  MUX2X1 _10575_ (
    .A( mem_backbone_0.pmem_dout_bckup_11_ ),
    .B(pmem_dout_11_),
    .S(_03925_),
    .Y(_03937_)
  );
  INVX1 _10576_ (
    .A(_03937_),
    .Y(_03731_)
  );
  MUX2X1 _10577_ (
    .A( mem_backbone_0.pmem_dout_bckup_12_ ),
    .B(pmem_dout_12_),
    .S(_03925_),
    .Y(_03938_)
  );
  INVX1 _10578_ (
    .A(_03938_),
    .Y(_03732_)
  );
  MUX2X1 _10579_ (
    .A( mem_backbone_0.pmem_dout_bckup_13_ ),
    .B(pmem_dout_13_),
    .S(_03925_),
    .Y(_03939_)
  );
  INVX1 _10580_ (
    .A(_03939_),
    .Y(_03733_)
  );
  MUX2X1 _10581_ (
    .A( mem_backbone_0.pmem_dout_bckup_14_ ),
    .B(pmem_dout_14_),
    .S(_03925_),
    .Y(_03940_)
  );
  INVX1 _10582_ (
    .A(_03940_),
    .Y(_03734_)
  );
  MUX2X1 _10583_ (
    .A( mem_backbone_0.pmem_dout_bckup_15_ ),
    .B(pmem_dout_15_),
    .S(_03925_),
    .Y(_03941_)
  );
  INVX1 _10584_ (
    .A(_03941_),
    .Y(_03735_)
  );
  NOR2X1 _10585_ (
    .A( mem_backbone_0.fe_pmem_en_dly ),
    .B(_03818_),
    .Y(_03942_)
  );
  NAND2X1 _10586_ (
    .A(_03737_),
    .B( mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_03943_)
  );
  OAI21X1 _10587_ (
    .A(_03942_),
    .B(_03943_),
    .C(_03925_),
    .Y(_03736_)
  );
  DFFSR _10588_ (
    .CLK(dco_clk),
    .D(_03720_),
    .Q( mem_backbone_0.pmem_dout_bckup_0_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10589_ (
    .CLK(dco_clk),
    .D(_03721_),
    .Q( mem_backbone_0.pmem_dout_bckup_1_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10590_ (
    .CLK(dco_clk),
    .D(_03722_),
    .Q( mem_backbone_0.pmem_dout_bckup_2_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10591_ (
    .CLK(dco_clk),
    .D(_03723_),
    .Q( mem_backbone_0.pmem_dout_bckup_3_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10592_ (
    .CLK(dco_clk),
    .D(_03724_),
    .Q( mem_backbone_0.pmem_dout_bckup_4_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10593_ (
    .CLK(dco_clk),
    .D(_03725_),
    .Q( mem_backbone_0.pmem_dout_bckup_5_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10594_ (
    .CLK(dco_clk),
    .D(_03726_),
    .Q( mem_backbone_0.pmem_dout_bckup_6_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10595_ (
    .CLK(dco_clk),
    .D(_03727_),
    .Q( mem_backbone_0.pmem_dout_bckup_7_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10596_ (
    .CLK(dco_clk),
    .D(_03728_),
    .Q( mem_backbone_0.pmem_dout_bckup_8_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10597_ (
    .CLK(dco_clk),
    .D(_03729_),
    .Q( mem_backbone_0.pmem_dout_bckup_9_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10598_ (
    .CLK(dco_clk),
    .D(_03730_),
    .Q( mem_backbone_0.pmem_dout_bckup_10_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10599_ (
    .CLK(dco_clk),
    .D(_03731_),
    .Q( mem_backbone_0.pmem_dout_bckup_11_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10600_ (
    .CLK(dco_clk),
    .D(_03732_),
    .Q( mem_backbone_0.pmem_dout_bckup_12_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10601_ (
    .CLK(dco_clk),
    .D(_03733_),
    .Q( mem_backbone_0.pmem_dout_bckup_13_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10602_ (
    .CLK(dco_clk),
    .D(_03734_),
    .Q( mem_backbone_0.pmem_dout_bckup_14_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10603_ (
    .CLK(dco_clk),
    .D(_03735_),
    .Q( mem_backbone_0.pmem_dout_bckup_15_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10604_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.ext_per_en ),
    .Q( mem_backbone_0.ext_mem_din_sel ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10605_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.ext_pmem_en ),
    .Q(_03718_),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10606_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.eu_per_en ),
    .Q( mem_backbone_0.eu_mdb_in_sel_0_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10607_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.eu_pmem_en ),
    .Q( mem_backbone_0.eu_mdb_in_sel_1_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10608_ (
    .CLK(dco_clk),
    .D(_03736_),
    .Q( mem_backbone_0.pmem_dout_bckup_sel ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10609_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.fe_pmem_en ),
    .Q( mem_backbone_0.fe_pmem_en_dly ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10610_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_0_ ),
    .Q( mem_backbone_0.per_dout_val_0_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10611_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_1_ ),
    .Q( mem_backbone_0.per_dout_val_1_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10612_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_2_ ),
    .Q( mem_backbone_0.per_dout_val_2_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10613_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_3_ ),
    .Q( mem_backbone_0.per_dout_val_3_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10614_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_4_ ),
    .Q( mem_backbone_0.per_dout_val_4_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10615_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_5_ ),
    .Q( mem_backbone_0.per_dout_val_5_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10616_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_6_ ),
    .Q( mem_backbone_0.per_dout_val_6_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10617_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_7_ ),
    .Q( mem_backbone_0.per_dout_val_7_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10618_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_8_ ),
    .Q( mem_backbone_0.per_dout_val_8_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10619_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_9_ ),
    .Q( mem_backbone_0.per_dout_val_9_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10620_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_10_ ),
    .Q( mem_backbone_0.per_dout_val_10_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10621_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_11_ ),
    .Q( mem_backbone_0.per_dout_val_11_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10622_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_12_ ),
    .Q( mem_backbone_0.per_dout_val_12_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10623_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_13_ ),
    .Q( mem_backbone_0.per_dout_val_13_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10624_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_14_ ),
    .Q( mem_backbone_0.per_dout_val_14_ ),
    .R(_03719_),
    .S(1'h1)
  );
  DFFSR _10625_ (
    .CLK(dco_clk),
    .D( mem_backbone_0.per_dout_15_ ),
    .Q( mem_backbone_0.per_dout_val_15_ ),
    .R(_03719_),
    .S(1'h1)
  );
  INVX1 _10626_ (
    .A( multiplier_0.cycle_1_ ),
    .Y(_04588_)
  );
  INVX1 _10627_ (
    .A( multiplier_0.cycle_0_ ),
    .Y(_04589_)
  );
  INVX1 _10628_ (
    .A(_05634_),
    .Y(_04590_)
  );
  INVX1 _10629_ (
    .A(_05637_),
    .Y(_04591_)
  );
  INVX1 _10630_ (
    .A(_05639_),
    .Y(_04592_)
  );
  INVX1 _10631_ (
    .A(_05640_),
    .Y(_04593_)
  );
  INVX1 _10632_ (
    .A(_05633_),
    .Y(_04594_)
  );
  INVX1 _10633_ (
    .A( multiplier_0.op2_0_ ),
    .Y(_04595_)
  );
  INVX1 _10634_ (
    .A( multiplier_0.op1_1_ ),
    .Y(_04596_)
  );
  INVX1 _10635_ (
    .A( multiplier_0.op2_1_ ),
    .Y(_04597_)
  );
  INVX1 _10636_ (
    .A( multiplier_0.reslo_2_ ),
    .Y(_04598_)
  );
  INVX1 _10637_ (
    .A( multiplier_0.op1_2_ ),
    .Y(_04599_)
  );
  INVX1 _10638_ (
    .A( multiplier_0.op2_2_ ),
    .Y(_04600_)
  );
  INVX1 _10639_ (
    .A( multiplier_0.op1_3_ ),
    .Y(_04601_)
  );
  INVX1 _10640_ (
    .A( multiplier_0.op2_3_ ),
    .Y(_04602_)
  );
  INVX1 _10641_ (
    .A( multiplier_0.op1_4_ ),
    .Y(_04603_)
  );
  INVX1 _10642_ (
    .A( multiplier_0.op2_4_ ),
    .Y(_04604_)
  );
  INVX1 _10643_ (
    .A( multiplier_0.op1_5_ ),
    .Y(_04605_)
  );
  INVX1 _10644_ (
    .A( multiplier_0.op2_5_ ),
    .Y(_04606_)
  );
  INVX1 _10645_ (
    .A( multiplier_0.op1_6_ ),
    .Y(_04607_)
  );
  INVX1 _10646_ (
    .A( multiplier_0.op2_6_ ),
    .Y(_04608_)
  );
  INVX1 _10647_ (
    .A( multiplier_0.op1_7_ ),
    .Y(_04609_)
  );
  INVX1 _10648_ (
    .A( multiplier_0.op2_7_ ),
    .Y(_04610_)
  );
  INVX1 _10649_ (
    .A( multiplier_0.op1_8_ ),
    .Y(_04611_)
  );
  INVX1 _10650_ (
    .A( multiplier_0.reslo_11_ ),
    .Y(_04612_)
  );
  INVX1 _10651_ (
    .A( multiplier_0.op1_14_ ),
    .Y(_04613_)
  );
  INVX1 _10652_ (
    .A( multiplier_0.reslo_15_ ),
    .Y(_04614_)
  );
  INVX1 _10653_ (
    .A( multiplier_0.reshi_3_ ),
    .Y(_04615_)
  );
  INVX1 _10654_ (
    .A( multiplier_0.reshi_5_ ),
    .Y(_04616_)
  );
  INVX1 _10655_ (
    .A( multiplier_0.reshi_7_ ),
    .Y(_04617_)
  );
  INVX1 _10656_ (
    .A( multiplier_0.reshi_15_ ),
    .Y(_04618_)
  );
  INVX1 _10657_ (
    .A( multiplier_0.sumext_0_ ),
    .Y(_04619_)
  );
  INVX1 _10658_ (
    .A(_05695_),
    .Y(_03944_)
  );
  NOR2X1 _10659_ (
    .A(_05661_),
    .B(_05660_),
    .Y(_04620_)
  );
  OR2X1 _10660_ (
    .A(_05632_),
    .B(1'h0),
    .Y(_04621_)
  );
  NAND2X1 _10661_ (
    .A(_04594_),
    .B(_05659_),
    .Y(_04622_)
  );
  NOR2X1 _10662_ (
    .A(_04621_),
    .B(_04622_),
    .Y(_04623_)
  );
  NOR2X1 _10663_ (
    .A(_05641_),
    .B(_04593_),
    .Y(_04624_)
  );
  NOR2X1 _10664_ (
    .A(_05631_),
    .B(_05642_),
    .Y(_04625_)
  );
  NAND2X1 _10665_ (
    .A(_04624_),
    .B(_04625_),
    .Y(_04626_)
  );
  NOR2X1 _10666_ (
    .A(_05639_),
    .B(_05638_),
    .Y(_04627_)
  );
  NAND3X1 _10667_ (
    .A(_05637_),
    .B(_05636_),
    .C(_04627_),
    .Y(_04628_)
  );
  NOR2X1 _10668_ (
    .A(_04626_),
    .B(_04628_),
    .Y(_04629_)
  );
  AND2X1 _10669_ (
    .A(_04623_),
    .B(_04629_),
    .Y(_04630_)
  );
  OAI21X1 _10670_ (
    .A(_05661_),
    .B(_05660_),
    .C(_04630_),
    .Y(_04631_)
  );
  NAND2X1 _10671_ (
    .A(_05635_),
    .B(_04590_),
    .Y(_04632_)
  );
  OR2X1 _10672_ (
    .A(_05630_),
    .B(_04632_),
    .Y(_04633_)
  );
  OR2X1 _10673_ (
    .A(_04631_),
    .B(_04633_),
    .Y(_04634_)
  );
  INVX1 _10674_ (
    .A(_04634_),
    .Y( multiplier_0.op2_wr )
  );
  NOR2X1 _10675_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.sign_sel ),
    .Y(_04635_)
  );
  NAND2X1 _10676_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_9_ ),
    .Y(_04636_)
  );
  MUX2X1 _10677_ (
    .A( multiplier_0.op2_9_ ),
    .B( multiplier_0.op2_1_ ),
    .S( multiplier_0.cycle_0_ ),
    .Y(_04637_)
  );
  OAI21X1 _10678_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04597_),
    .C(_04636_),
    .Y(_04638_)
  );
  NAND2X1 _10679_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_8_ ),
    .Y(_04639_)
  );
  NOR2X1 _10680_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04595_),
    .Y(_04640_)
  );
  MUX2X1 _10681_ (
    .A( multiplier_0.op2_8_ ),
    .B( multiplier_0.op2_0_ ),
    .S( multiplier_0.cycle_0_ ),
    .Y(_04641_)
  );
  OAI21X1 _10682_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04595_),
    .C(_04639_),
    .Y(_04642_)
  );
  AND2X1 _10683_ (
    .A( multiplier_0.sign_sel ),
    .B( multiplier_0.op1_15_ ),
    .Y(_04643_)
  );
  NAND2X1 _10684_ (
    .A( multiplier_0.sign_sel ),
    .B( multiplier_0.op1_15_ ),
    .Y(_04644_)
  );
  NAND2X1 _10685_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04642_),
    .Y(_04645_)
  );
  NOR2X1 _10686_ (
    .A(_04641_),
    .B(_04644_),
    .Y(_04646_)
  );
  NAND2X1 _10687_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04638_),
    .Y(_04647_)
  );
  INVX1 _10688_ (
    .A(_04647_),
    .Y(_04648_)
  );
  NAND2X1 _10689_ (
    .A(_04638_),
    .B(_04646_),
    .Y(_04649_)
  );
  NAND2X1 _10690_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_10_ ),
    .Y(_04650_)
  );
  OAI21X1 _10691_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04600_),
    .C(_04650_),
    .Y(_04651_)
  );
  NAND2X1 _10692_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04651_),
    .Y(_04652_)
  );
  NAND2X1 _10693_ (
    .A(_04643_),
    .B(_04651_),
    .Y(_04653_)
  );
  NOR2X1 _10694_ (
    .A(_04649_),
    .B(_04653_),
    .Y(_04654_)
  );
  OR2X1 _10695_ (
    .A(_04649_),
    .B(_04653_),
    .Y(_04655_)
  );
  NAND2X1 _10696_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_13_ ),
    .Y(_04656_)
  );
  OAI21X1 _10697_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04606_),
    .C(_04656_),
    .Y(_04657_)
  );
  NAND2X1 _10698_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04657_),
    .Y(_04658_)
  );
  NAND2X1 _10699_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_12_ ),
    .Y(_04659_)
  );
  OAI21X1 _10700_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04604_),
    .C(_04659_),
    .Y(_04660_)
  );
  NAND2X1 _10701_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04660_),
    .Y(_04661_)
  );
  NAND2X1 _10702_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_11_ ),
    .Y(_04662_)
  );
  OAI21X1 _10703_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04602_),
    .C(_04662_),
    .Y(_04663_)
  );
  NAND2X1 _10704_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04663_),
    .Y(_04664_)
  );
  NAND2X1 _10705_ (
    .A(_04643_),
    .B(_04663_),
    .Y(_04665_)
  );
  OR2X1 _10706_ (
    .A(_04661_),
    .B(_04665_),
    .Y(_04666_)
  );
  XNOR2X1 _10707_ (
    .A(_04661_),
    .B(_04665_),
    .Y(_04667_)
  );
  NAND2X1 _10708_ (
    .A(_04658_),
    .B(_04667_),
    .Y(_04668_)
  );
  OR2X1 _10709_ (
    .A(_04658_),
    .B(_04667_),
    .Y(_04669_)
  );
  NAND2X1 _10710_ (
    .A(_04668_),
    .B(_04669_),
    .Y(_04670_)
  );
  AOI21X1 _10711_ (
    .A(_04637_),
    .B(_04641_),
    .C(_04644_),
    .Y(_04671_)
  );
  AOI21X1 _10712_ (
    .A(_04643_),
    .B(_04651_),
    .C(_04671_),
    .Y(_04672_)
  );
  NOR2X1 _10713_ (
    .A(_04654_),
    .B(_04672_),
    .Y(_04673_)
  );
  NAND3X1 _10714_ (
    .A(_04668_),
    .B(_04669_),
    .C(_04673_),
    .Y(_04674_)
  );
  AND2X1 _10715_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04657_),
    .Y(_04675_)
  );
  NAND2X1 _10716_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04657_),
    .Y(_04676_)
  );
  OAI21X1 _10717_ (
    .A(_04660_),
    .B(_04663_),
    .C(_04643_),
    .Y(_04677_)
  );
  INVX1 _10718_ (
    .A(_04677_),
    .Y(_04678_)
  );
  OAI21X1 _10719_ (
    .A(_04661_),
    .B(_04665_),
    .C(_04678_),
    .Y(_04679_)
  );
  XNOR2X1 _10720_ (
    .A(_04675_),
    .B(_04679_),
    .Y(_04680_)
  );
  XNOR2X1 _10721_ (
    .A(_04673_),
    .B(_04680_),
    .Y(_04681_)
  );
  AOI21X1 _10722_ (
    .A(_04655_),
    .B(_04674_),
    .C(_04681_),
    .Y(_04682_)
  );
  INVX1 _10723_ (
    .A(_04682_),
    .Y(_04683_)
  );
  NAND2X1 _10724_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_15_ ),
    .Y(_04684_)
  );
  OAI21X1 _10725_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04610_),
    .C(_04684_),
    .Y(_04685_)
  );
  NAND2X1 _10726_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04685_),
    .Y(_04686_)
  );
  NAND2X1 _10727_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_14_ ),
    .Y(_04687_)
  );
  OAI21X1 _10728_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04608_),
    .C(_04687_),
    .Y(_04688_)
  );
  NAND2X1 _10729_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04688_),
    .Y(_04689_)
  );
  NAND2X1 _10730_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04685_),
    .Y(_04690_)
  );
  NAND2X1 _10731_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04688_),
    .Y(_04691_)
  );
  OR2X1 _10732_ (
    .A(_04686_),
    .B(_04689_),
    .Y(_04692_)
  );
  NAND3X1 _10733_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.op2_15_ ),
    .C( multiplier_0.sign_sel ),
    .Y(_04693_)
  );
  NOR2X1 _10734_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04693_),
    .Y(_04694_)
  );
  NAND2X1 _10735_ (
    .A(_04686_),
    .B(_04689_),
    .Y(_04695_)
  );
  OAI21X1 _10736_ (
    .A(_04690_),
    .B(_04691_),
    .C(_04695_),
    .Y(_04696_)
  );
  NAND3X1 _10737_ (
    .A(_04692_),
    .B(_04694_),
    .C(_04695_),
    .Y(_04697_)
  );
  OAI21X1 _10738_ (
    .A(_04690_),
    .B(_04691_),
    .C(_04697_),
    .Y(_04698_)
  );
  OR2X1 _10739_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04693_),
    .Y(_04699_)
  );
  NAND2X1 _10740_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04688_),
    .Y(_04700_)
  );
  NAND2X1 _10741_ (
    .A(_04690_),
    .B(_04700_),
    .Y(_04701_)
  );
  NAND2X1 _10742_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04685_),
    .Y(_04702_)
  );
  OAI21X1 _10743_ (
    .A(_04689_),
    .B(_04702_),
    .C(_04701_),
    .Y(_04703_)
  );
  OAI21X1 _10744_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04693_),
    .C(_04703_),
    .Y(_04704_)
  );
  OR2X1 _10745_ (
    .A(_04699_),
    .B(_04703_),
    .Y(_04705_)
  );
  NAND2X1 _10746_ (
    .A(_04704_),
    .B(_04705_),
    .Y(_04706_)
  );
  AND2X1 _10747_ (
    .A(_04666_),
    .B(_04669_),
    .Y(_04707_)
  );
  NOR2X1 _10748_ (
    .A(_04706_),
    .B(_04707_),
    .Y(_04708_)
  );
  XNOR2X1 _10749_ (
    .A(_04706_),
    .B(_04707_),
    .Y(_04709_)
  );
  AOI21X1 _10750_ (
    .A(_04692_),
    .B(_04697_),
    .C(_04709_),
    .Y(_04710_)
  );
  XOR2X1 _10751_ (
    .A(_04698_),
    .B(_04709_),
    .Y(_04711_)
  );
  NAND3X1 _10752_ (
    .A(_04655_),
    .B(_04674_),
    .C(_04681_),
    .Y(_04712_)
  );
  NAND2X1 _10753_ (
    .A(_04683_),
    .B(_04712_),
    .Y(_04713_)
  );
  OAI21X1 _10754_ (
    .A(_04711_),
    .B(_04713_),
    .C(_04683_),
    .Y(_04714_)
  );
  OAI21X1 _10755_ (
    .A(_04689_),
    .B(_04702_),
    .C(_04705_),
    .Y(_04715_)
  );
  OR2X1 _10756_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04693_),
    .Y(_04716_)
  );
  NAND2X1 _10757_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04688_),
    .Y(_04717_)
  );
  NAND2X1 _10758_ (
    .A(_04702_),
    .B(_04717_),
    .Y(_04718_)
  );
  NAND2X1 _10759_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04685_),
    .Y(_04719_)
  );
  OAI21X1 _10760_ (
    .A(_04700_),
    .B(_04719_),
    .C(_04718_),
    .Y(_04720_)
  );
  OAI21X1 _10761_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04693_),
    .C(_04720_),
    .Y(_04721_)
  );
  OR2X1 _10762_ (
    .A(_04716_),
    .B(_04720_),
    .Y(_04722_)
  );
  NAND2X1 _10763_ (
    .A(_04721_),
    .B(_04722_),
    .Y(_04723_)
  );
  OAI21X1 _10764_ (
    .A(_04676_),
    .B(_04677_),
    .C(_04666_),
    .Y(_04724_)
  );
  INVX1 _10765_ (
    .A(_04724_),
    .Y(_04725_)
  );
  NOR2X1 _10766_ (
    .A(_04723_),
    .B(_04725_),
    .Y(_04726_)
  );
  NAND2X1 _10767_ (
    .A(_04723_),
    .B(_04725_),
    .Y(_04727_)
  );
  XNOR2X1 _10768_ (
    .A(_04723_),
    .B(_04724_),
    .Y(_04728_)
  );
  XNOR2X1 _10769_ (
    .A(_04715_),
    .B(_04728_),
    .Y(_04729_)
  );
  NAND2X1 _10770_ (
    .A(_04643_),
    .B(_04657_),
    .Y(_04730_)
  );
  MUX2X1 _10771_ (
    .A(_04730_),
    .B(_04675_),
    .S(_04679_),
    .Y(_04731_)
  );
  NAND2X1 _10772_ (
    .A(_04654_),
    .B(_04731_),
    .Y(_04732_)
  );
  MUX2X1 _10773_ (
    .A(_04654_),
    .B(_04672_),
    .S(_04731_),
    .Y(_04733_)
  );
  INVX1 _10774_ (
    .A(_04733_),
    .Y(_04734_)
  );
  NOR2X1 _10775_ (
    .A(_04729_),
    .B(_04734_),
    .Y(_04735_)
  );
  XNOR2X1 _10776_ (
    .A(_04729_),
    .B(_04733_),
    .Y(_04736_)
  );
  NAND2X1 _10777_ (
    .A(_04714_),
    .B(_04736_),
    .Y(_04737_)
  );
  NOR2X1 _10778_ (
    .A(_04708_),
    .B(_04710_),
    .Y(_04738_)
  );
  XNOR2X1 _10779_ (
    .A(_04714_),
    .B(_04736_),
    .Y(_04739_)
  );
  OAI21X1 _10780_ (
    .A(_04738_),
    .B(_04739_),
    .C(_04737_),
    .Y(_04740_)
  );
  AOI21X1 _10781_ (
    .A(_04715_),
    .B(_04727_),
    .C(_04726_),
    .Y(_04741_)
  );
  AOI21X1 _10782_ (
    .A(_04654_),
    .B(_04731_),
    .C(_04735_),
    .Y(_04742_)
  );
  OAI21X1 _10783_ (
    .A(_04700_),
    .B(_04719_),
    .C(_04722_),
    .Y(_04743_)
  );
  OR2X1 _10784_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04693_),
    .Y(_04744_)
  );
  NAND2X1 _10785_ (
    .A(_04643_),
    .B(_04688_),
    .Y(_04745_)
  );
  NAND2X1 _10786_ (
    .A(_04719_),
    .B(_04745_),
    .Y(_04746_)
  );
  OR2X1 _10787_ (
    .A(_04719_),
    .B(_04745_),
    .Y(_04747_)
  );
  NAND2X1 _10788_ (
    .A(_04746_),
    .B(_04747_),
    .Y(_04748_)
  );
  NOR2X1 _10789_ (
    .A(_04744_),
    .B(_04748_),
    .Y(_04749_)
  );
  XNOR2X1 _10790_ (
    .A(_04744_),
    .B(_04748_),
    .Y(_04750_)
  );
  XNOR2X1 _10791_ (
    .A(_04724_),
    .B(_04750_),
    .Y(_04751_)
  );
  NAND2X1 _10792_ (
    .A(_04743_),
    .B(_04751_),
    .Y(_04752_)
  );
  XNOR2X1 _10793_ (
    .A(_04743_),
    .B(_04751_),
    .Y(_04753_)
  );
  XNOR2X1 _10794_ (
    .A(_04734_),
    .B(_04753_),
    .Y(_04754_)
  );
  XNOR2X1 _10795_ (
    .A(_04742_),
    .B(_04754_),
    .Y(_04755_)
  );
  OR2X1 _10796_ (
    .A(_04741_),
    .B(_04755_),
    .Y(_04756_)
  );
  XOR2X1 _10797_ (
    .A(_04741_),
    .B(_04755_),
    .Y(_04757_)
  );
  NAND2X1 _10798_ (
    .A(_04740_),
    .B(_04757_),
    .Y(_04758_)
  );
  XNOR2X1 _10799_ (
    .A(_04740_),
    .B(_04757_),
    .Y(_04759_)
  );
  XOR2X1 _10800_ (
    .A(_04738_),
    .B(_04739_),
    .Y(_04760_)
  );
  NAND2X1 _10801_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04657_),
    .Y(_04761_)
  );
  NAND2X1 _10802_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04660_),
    .Y(_04762_)
  );
  NAND2X1 _10803_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04663_),
    .Y(_04763_)
  );
  XNOR2X1 _10804_ (
    .A(_04664_),
    .B(_04762_),
    .Y(_04764_)
  );
  XNOR2X1 _10805_ (
    .A(_04761_),
    .B(_04764_),
    .Y(_04765_)
  );
  OAI21X1 _10806_ (
    .A(_04672_),
    .B(_04765_),
    .C(_04655_),
    .Y(_04766_)
  );
  OAI21X1 _10807_ (
    .A(_04654_),
    .B(_04672_),
    .C(_04670_),
    .Y(_04767_)
  );
  AND2X1 _10808_ (
    .A(_04674_),
    .B(_04767_),
    .Y(_04768_)
  );
  NAND2X1 _10809_ (
    .A(_04766_),
    .B(_04768_),
    .Y(_04769_)
  );
  NAND2X1 _10810_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04685_),
    .Y(_04770_)
  );
  NAND2X1 _10811_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04688_),
    .Y(_04771_)
  );
  OR2X1 _10812_ (
    .A(_04691_),
    .B(_04770_),
    .Y(_04772_)
  );
  NOR2X1 _10813_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04693_),
    .Y(_04773_)
  );
  INVX1 _10814_ (
    .A(_04773_),
    .Y(_04774_)
  );
  NAND2X1 _10815_ (
    .A(_04691_),
    .B(_04770_),
    .Y(_04775_)
  );
  OAI21X1 _10816_ (
    .A(_04686_),
    .B(_04771_),
    .C(_04775_),
    .Y(_04776_)
  );
  OAI21X1 _10817_ (
    .A(_04774_),
    .B(_04776_),
    .C(_04772_),
    .Y(_04777_)
  );
  OAI21X1 _10818_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04693_),
    .C(_04696_),
    .Y(_04778_)
  );
  NAND2X1 _10819_ (
    .A(_04697_),
    .B(_04778_),
    .Y(_04779_)
  );
  OAI22X1 _10820_ (
    .A(_04661_),
    .B(_04763_),
    .C(_04764_),
    .D(_04761_),
    .Y(_04780_)
  );
  INVX1 _10821_ (
    .A(_04780_),
    .Y(_04781_)
  );
  XNOR2X1 _10822_ (
    .A(_04779_),
    .B(_04781_),
    .Y(_04782_)
  );
  INVX1 _10823_ (
    .A(_04782_),
    .Y(_04783_)
  );
  NAND2X1 _10824_ (
    .A(_04777_),
    .B(_04783_),
    .Y(_04784_)
  );
  XOR2X1 _10825_ (
    .A(_04777_),
    .B(_04782_),
    .Y(_04785_)
  );
  XNOR2X1 _10826_ (
    .A(_04766_),
    .B(_04768_),
    .Y(_04786_)
  );
  OAI21X1 _10827_ (
    .A(_04785_),
    .B(_04786_),
    .C(_04769_),
    .Y(_04787_)
  );
  XOR2X1 _10828_ (
    .A(_04711_),
    .B(_04713_),
    .Y(_04788_)
  );
  NAND2X1 _10829_ (
    .A(_04787_),
    .B(_04788_),
    .Y(_04789_)
  );
  OAI21X1 _10830_ (
    .A(_04779_),
    .B(_04781_),
    .C(_04784_),
    .Y(_04790_)
  );
  INVX1 _10831_ (
    .A(_04790_),
    .Y(_04791_)
  );
  XNOR2X1 _10832_ (
    .A(_04787_),
    .B(_04788_),
    .Y(_04792_)
  );
  OAI21X1 _10833_ (
    .A(_04791_),
    .B(_04792_),
    .C(_04789_),
    .Y(_04793_)
  );
  NAND2X1 _10834_ (
    .A(_04760_),
    .B(_04793_),
    .Y(_04794_)
  );
  NOR2X1 _10835_ (
    .A(_04759_),
    .B(_04794_),
    .Y(_04795_)
  );
  XOR2X1 _10836_ (
    .A(_04760_),
    .B(_04793_),
    .Y(_04796_)
  );
  XNOR2X1 _10837_ (
    .A(_04790_),
    .B(_04792_),
    .Y(_04797_)
  );
  NAND2X1 _10838_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04651_),
    .Y(_04798_)
  );
  OAI21X1 _10839_ (
    .A(_04646_),
    .B(_04648_),
    .C(_04649_),
    .Y(_04799_)
  );
  OAI21X1 _10840_ (
    .A(_04798_),
    .B(_04799_),
    .C(_04649_),
    .Y(_04800_)
  );
  NAND2X1 _10841_ (
    .A(_04649_),
    .B(_04671_),
    .Y(_04801_)
  );
  NAND2X1 _10842_ (
    .A(_04652_),
    .B(_04801_),
    .Y(_04802_)
  );
  OAI21X1 _10843_ (
    .A(_04653_),
    .B(_04801_),
    .C(_04802_),
    .Y(_04803_)
  );
  INVX1 _10844_ (
    .A(_04803_),
    .Y(_04804_)
  );
  NAND2X1 _10845_ (
    .A(_04800_),
    .B(_04804_),
    .Y(_04805_)
  );
  NAND2X1 _10846_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04657_),
    .Y(_04806_)
  );
  NAND2X1 _10847_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04660_),
    .Y(_04807_)
  );
  NAND2X1 _10848_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04663_),
    .Y(_04808_)
  );
  XNOR2X1 _10849_ (
    .A(_04763_),
    .B(_04807_),
    .Y(_04809_)
  );
  XOR2X1 _10850_ (
    .A(_04806_),
    .B(_04809_),
    .Y(_04810_)
  );
  XNOR2X1 _10851_ (
    .A(_04800_),
    .B(_04803_),
    .Y(_04811_)
  );
  NAND2X1 _10852_ (
    .A(_04810_),
    .B(_04811_),
    .Y(_04812_)
  );
  XOR2X1 _10853_ (
    .A(_04673_),
    .B(_04765_),
    .Y(_04813_)
  );
  AOI21X1 _10854_ (
    .A(_04805_),
    .B(_04812_),
    .C(_04813_),
    .Y(_04814_)
  );
  INVX1 _10855_ (
    .A(_04814_),
    .Y(_04815_)
  );
  NAND2X1 _10856_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04685_),
    .Y(_04816_)
  );
  NAND2X1 _10857_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04688_),
    .Y(_04817_)
  );
  NOR2X1 _10858_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04693_),
    .Y(_04818_)
  );
  INVX1 _10859_ (
    .A(_04818_),
    .Y(_04819_)
  );
  NAND2X1 _10860_ (
    .A(_04771_),
    .B(_04816_),
    .Y(_04820_)
  );
  OAI21X1 _10861_ (
    .A(_04770_),
    .B(_04817_),
    .C(_04820_),
    .Y(_04821_)
  );
  OAI22X1 _10862_ (
    .A(_04770_),
    .B(_04817_),
    .C(_04819_),
    .D(_04821_),
    .Y(_04822_)
  );
  XNOR2X1 _10863_ (
    .A(_04774_),
    .B(_04776_),
    .Y(_04823_)
  );
  OAI22X1 _10864_ (
    .A(_04762_),
    .B(_04808_),
    .C(_04809_),
    .D(_04806_),
    .Y(_04824_)
  );
  INVX1 _10865_ (
    .A(_04824_),
    .Y(_04825_)
  );
  XNOR2X1 _10866_ (
    .A(_04823_),
    .B(_04825_),
    .Y(_04826_)
  );
  INVX1 _10867_ (
    .A(_04826_),
    .Y(_04827_)
  );
  NAND2X1 _10868_ (
    .A(_04822_),
    .B(_04827_),
    .Y(_04828_)
  );
  XOR2X1 _10869_ (
    .A(_04822_),
    .B(_04826_),
    .Y(_04829_)
  );
  NAND3X1 _10870_ (
    .A(_04805_),
    .B(_04812_),
    .C(_04813_),
    .Y(_04830_)
  );
  NAND2X1 _10871_ (
    .A(_04815_),
    .B(_04830_),
    .Y(_04831_)
  );
  OAI21X1 _10872_ (
    .A(_04829_),
    .B(_04831_),
    .C(_04815_),
    .Y(_04832_)
  );
  XOR2X1 _10873_ (
    .A(_04785_),
    .B(_04786_),
    .Y(_04833_)
  );
  NAND2X1 _10874_ (
    .A(_04832_),
    .B(_04833_),
    .Y(_04834_)
  );
  OAI21X1 _10875_ (
    .A(_04823_),
    .B(_04825_),
    .C(_04828_),
    .Y(_04835_)
  );
  INVX1 _10876_ (
    .A(_04835_),
    .Y(_04836_)
  );
  XNOR2X1 _10877_ (
    .A(_04832_),
    .B(_04833_),
    .Y(_04837_)
  );
  OAI21X1 _10878_ (
    .A(_04836_),
    .B(_04837_),
    .C(_04834_),
    .Y(_04838_)
  );
  NAND2X1 _10879_ (
    .A(_04797_),
    .B(_04838_),
    .Y(_04839_)
  );
  NAND3X1 _10880_ (
    .A(_04796_),
    .B(_04797_),
    .C(_04838_),
    .Y(_04840_)
  );
  XNOR2X1 _10881_ (
    .A(_04796_),
    .B(_04839_),
    .Y(_04841_)
  );
  INVX1 _10882_ (
    .A(_04841_),
    .Y(_04842_)
  );
  XNOR2X1 _10883_ (
    .A(_04797_),
    .B(_04838_),
    .Y(_04843_)
  );
  XNOR2X1 _10884_ (
    .A(_04835_),
    .B(_04837_),
    .Y(_04844_)
  );
  NAND2X1 _10885_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04642_),
    .Y(_04845_)
  );
  NAND2X1 _10886_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04651_),
    .Y(_04846_)
  );
  OAI21X1 _10887_ (
    .A(_04613_),
    .B(_04637_),
    .C(_04645_),
    .Y(_04847_)
  );
  OAI21X1 _10888_ (
    .A(_04647_),
    .B(_04845_),
    .C(_04847_),
    .Y(_04848_)
  );
  OAI22X1 _10889_ (
    .A(_04647_),
    .B(_04845_),
    .C(_04846_),
    .D(_04848_),
    .Y(_04849_)
  );
  XNOR2X1 _10890_ (
    .A(_04798_),
    .B(_04799_),
    .Y(_04850_)
  );
  INVX1 _10891_ (
    .A(_04850_),
    .Y(_04851_)
  );
  NAND2X1 _10892_ (
    .A(_04849_),
    .B(_04851_),
    .Y(_04852_)
  );
  NAND2X1 _10893_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04657_),
    .Y(_04853_)
  );
  NAND2X1 _10894_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04660_),
    .Y(_04854_)
  );
  NAND2X1 _10895_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04663_),
    .Y(_04855_)
  );
  XNOR2X1 _10896_ (
    .A(_04808_),
    .B(_04854_),
    .Y(_04856_)
  );
  XNOR2X1 _10897_ (
    .A(_04853_),
    .B(_04856_),
    .Y(_04857_)
  );
  XOR2X1 _10898_ (
    .A(_04849_),
    .B(_04850_),
    .Y(_04858_)
  );
  OAI21X1 _10899_ (
    .A(_04857_),
    .B(_04858_),
    .C(_04852_),
    .Y(_04859_)
  );
  XOR2X1 _10900_ (
    .A(_04810_),
    .B(_04811_),
    .Y(_04860_)
  );
  NAND2X1 _10901_ (
    .A(_04859_),
    .B(_04860_),
    .Y(_04861_)
  );
  NAND2X1 _10902_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04685_),
    .Y(_04862_)
  );
  NAND2X1 _10903_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04688_),
    .Y(_04863_)
  );
  NOR2X1 _10904_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04693_),
    .Y(_04864_)
  );
  INVX1 _10905_ (
    .A(_04864_),
    .Y(_04865_)
  );
  NAND2X1 _10906_ (
    .A(_04817_),
    .B(_04862_),
    .Y(_04866_)
  );
  OAI21X1 _10907_ (
    .A(_04816_),
    .B(_04863_),
    .C(_04866_),
    .Y(_04867_)
  );
  OAI22X1 _10908_ (
    .A(_04816_),
    .B(_04863_),
    .C(_04865_),
    .D(_04867_),
    .Y(_04868_)
  );
  XNOR2X1 _10909_ (
    .A(_04819_),
    .B(_04821_),
    .Y(_04869_)
  );
  OAI22X1 _10910_ (
    .A(_04807_),
    .B(_04855_),
    .C(_04856_),
    .D(_04853_),
    .Y(_04870_)
  );
  INVX1 _10911_ (
    .A(_04870_),
    .Y(_04871_)
  );
  XOR2X1 _10912_ (
    .A(_04869_),
    .B(_04870_),
    .Y(_04872_)
  );
  INVX1 _10913_ (
    .A(_04872_),
    .Y(_04873_)
  );
  NAND2X1 _10914_ (
    .A(_04868_),
    .B(_04873_),
    .Y(_04874_)
  );
  XOR2X1 _10915_ (
    .A(_04868_),
    .B(_04872_),
    .Y(_04875_)
  );
  XNOR2X1 _10916_ (
    .A(_04859_),
    .B(_04860_),
    .Y(_04876_)
  );
  OAI21X1 _10917_ (
    .A(_04875_),
    .B(_04876_),
    .C(_04861_),
    .Y(_04877_)
  );
  XOR2X1 _10918_ (
    .A(_04829_),
    .B(_04831_),
    .Y(_04878_)
  );
  NAND2X1 _10919_ (
    .A(_04877_),
    .B(_04878_),
    .Y(_04879_)
  );
  OAI21X1 _10920_ (
    .A(_04869_),
    .B(_04871_),
    .C(_04874_),
    .Y(_04880_)
  );
  INVX1 _10921_ (
    .A(_04880_),
    .Y(_04881_)
  );
  XNOR2X1 _10922_ (
    .A(_04877_),
    .B(_04878_),
    .Y(_04882_)
  );
  OAI21X1 _10923_ (
    .A(_04881_),
    .B(_04882_),
    .C(_04879_),
    .Y(_04883_)
  );
  NAND2X1 _10924_ (
    .A(_04844_),
    .B(_04883_),
    .Y(_04884_)
  );
  NOR2X1 _10925_ (
    .A(_04843_),
    .B(_04884_),
    .Y(_04885_)
  );
  XOR2X1 _10926_ (
    .A(_04843_),
    .B(_04884_),
    .Y(_04886_)
  );
  XNOR2X1 _10927_ (
    .A(_04844_),
    .B(_04883_),
    .Y(_04887_)
  );
  XNOR2X1 _10928_ (
    .A(_04880_),
    .B(_04882_),
    .Y(_04888_)
  );
  NAND2X1 _10929_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04638_),
    .Y(_04889_)
  );
  NAND2X1 _10930_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04642_),
    .Y(_04890_)
  );
  NAND2X1 _10931_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04651_),
    .Y(_04891_)
  );
  XNOR2X1 _10932_ (
    .A(_04845_),
    .B(_04889_),
    .Y(_04892_)
  );
  OR2X1 _10933_ (
    .A(_04891_),
    .B(_04892_),
    .Y(_04893_)
  );
  OAI21X1 _10934_ (
    .A(_04845_),
    .B(_04889_),
    .C(_04893_),
    .Y(_04894_)
  );
  XNOR2X1 _10935_ (
    .A(_04846_),
    .B(_04848_),
    .Y(_04895_)
  );
  INVX1 _10936_ (
    .A(_04895_),
    .Y(_04896_)
  );
  NAND2X1 _10937_ (
    .A(_04894_),
    .B(_04896_),
    .Y(_04897_)
  );
  NAND2X1 _10938_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04657_),
    .Y(_04898_)
  );
  NAND2X1 _10939_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04660_),
    .Y(_04899_)
  );
  NAND2X1 _10940_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04663_),
    .Y(_04900_)
  );
  XNOR2X1 _10941_ (
    .A(_04855_),
    .B(_04899_),
    .Y(_04901_)
  );
  XNOR2X1 _10942_ (
    .A(_04898_),
    .B(_04901_),
    .Y(_04902_)
  );
  XOR2X1 _10943_ (
    .A(_04894_),
    .B(_04895_),
    .Y(_04903_)
  );
  OAI21X1 _10944_ (
    .A(_04902_),
    .B(_04903_),
    .C(_04897_),
    .Y(_04904_)
  );
  XOR2X1 _10945_ (
    .A(_04857_),
    .B(_04858_),
    .Y(_04905_)
  );
  NAND2X1 _10946_ (
    .A(_04904_),
    .B(_04905_),
    .Y(_04906_)
  );
  NAND2X1 _10947_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04685_),
    .Y(_04907_)
  );
  NAND2X1 _10948_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04688_),
    .Y(_04908_)
  );
  NOR2X1 _10949_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04693_),
    .Y(_04909_)
  );
  INVX1 _10950_ (
    .A(_04909_),
    .Y(_04910_)
  );
  NAND2X1 _10951_ (
    .A(_04863_),
    .B(_04907_),
    .Y(_04911_)
  );
  OAI21X1 _10952_ (
    .A(_04862_),
    .B(_04908_),
    .C(_04911_),
    .Y(_04912_)
  );
  OAI22X1 _10953_ (
    .A(_04862_),
    .B(_04908_),
    .C(_04910_),
    .D(_04912_),
    .Y(_04913_)
  );
  XNOR2X1 _10954_ (
    .A(_04865_),
    .B(_04867_),
    .Y(_04914_)
  );
  OAI22X1 _10955_ (
    .A(_04854_),
    .B(_04900_),
    .C(_04901_),
    .D(_04898_),
    .Y(_04915_)
  );
  INVX1 _10956_ (
    .A(_04915_),
    .Y(_04916_)
  );
  XNOR2X1 _10957_ (
    .A(_04914_),
    .B(_04916_),
    .Y(_04917_)
  );
  INVX1 _10958_ (
    .A(_04917_),
    .Y(_04918_)
  );
  NAND2X1 _10959_ (
    .A(_04913_),
    .B(_04918_),
    .Y(_04919_)
  );
  XOR2X1 _10960_ (
    .A(_04913_),
    .B(_04917_),
    .Y(_04920_)
  );
  XNOR2X1 _10961_ (
    .A(_04904_),
    .B(_04905_),
    .Y(_04921_)
  );
  OAI21X1 _10962_ (
    .A(_04920_),
    .B(_04921_),
    .C(_04906_),
    .Y(_04922_)
  );
  XOR2X1 _10963_ (
    .A(_04875_),
    .B(_04876_),
    .Y(_04923_)
  );
  NAND2X1 _10964_ (
    .A(_04922_),
    .B(_04923_),
    .Y(_04924_)
  );
  OAI21X1 _10965_ (
    .A(_04914_),
    .B(_04916_),
    .C(_04919_),
    .Y(_04925_)
  );
  INVX1 _10966_ (
    .A(_04925_),
    .Y(_04926_)
  );
  XNOR2X1 _10967_ (
    .A(_04922_),
    .B(_04923_),
    .Y(_04927_)
  );
  OAI21X1 _10968_ (
    .A(_04926_),
    .B(_04927_),
    .C(_04924_),
    .Y(_04928_)
  );
  NAND2X1 _10969_ (
    .A(_04888_),
    .B(_04928_),
    .Y(_04929_)
  );
  OR2X1 _10970_ (
    .A(_04887_),
    .B(_04929_),
    .Y(_04930_)
  );
  XOR2X1 _10971_ (
    .A(_04887_),
    .B(_04929_),
    .Y(_04931_)
  );
  INVX1 _10972_ (
    .A(_04931_),
    .Y(_04932_)
  );
  XNOR2X1 _10973_ (
    .A(_04888_),
    .B(_04928_),
    .Y(_04933_)
  );
  XNOR2X1 _10974_ (
    .A(_04925_),
    .B(_04927_),
    .Y(_04934_)
  );
  NAND2X1 _10975_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04638_),
    .Y(_04935_)
  );
  NAND2X1 _10976_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04642_),
    .Y(_04936_)
  );
  NAND2X1 _10977_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04651_),
    .Y(_04937_)
  );
  XNOR2X1 _10978_ (
    .A(_04890_),
    .B(_04935_),
    .Y(_04938_)
  );
  OAI22X1 _10979_ (
    .A(_04889_),
    .B(_04936_),
    .C(_04937_),
    .D(_04938_),
    .Y(_04939_)
  );
  NAND2X1 _10980_ (
    .A(_04891_),
    .B(_04892_),
    .Y(_04940_)
  );
  NAND2X1 _10981_ (
    .A(_04893_),
    .B(_04940_),
    .Y(_04941_)
  );
  NAND3X1 _10982_ (
    .A(_04893_),
    .B(_04939_),
    .C(_04940_),
    .Y(_04942_)
  );
  NAND2X1 _10983_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04657_),
    .Y(_04943_)
  );
  NAND2X1 _10984_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04660_),
    .Y(_04944_)
  );
  NAND2X1 _10985_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04663_),
    .Y(_04945_)
  );
  XNOR2X1 _10986_ (
    .A(_04900_),
    .B(_04944_),
    .Y(_04946_)
  );
  XNOR2X1 _10987_ (
    .A(_04943_),
    .B(_04946_),
    .Y(_04947_)
  );
  XOR2X1 _10988_ (
    .A(_04939_),
    .B(_04941_),
    .Y(_04948_)
  );
  OAI21X1 _10989_ (
    .A(_04947_),
    .B(_04948_),
    .C(_04942_),
    .Y(_04949_)
  );
  XOR2X1 _10990_ (
    .A(_04902_),
    .B(_04903_),
    .Y(_04950_)
  );
  NAND2X1 _10991_ (
    .A(_04949_),
    .B(_04950_),
    .Y(_04951_)
  );
  NAND2X1 _10992_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04685_),
    .Y(_04952_)
  );
  NAND2X1 _10993_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04688_),
    .Y(_04953_)
  );
  NOR2X1 _10994_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04693_),
    .Y(_04954_)
  );
  INVX1 _10995_ (
    .A(_04954_),
    .Y(_04955_)
  );
  NAND2X1 _10996_ (
    .A(_04908_),
    .B(_04952_),
    .Y(_04956_)
  );
  OAI21X1 _10997_ (
    .A(_04907_),
    .B(_04953_),
    .C(_04956_),
    .Y(_04957_)
  );
  OAI22X1 _10998_ (
    .A(_04907_),
    .B(_04953_),
    .C(_04955_),
    .D(_04957_),
    .Y(_04958_)
  );
  XNOR2X1 _10999_ (
    .A(_04910_),
    .B(_04912_),
    .Y(_04959_)
  );
  OAI22X1 _11000_ (
    .A(_04899_),
    .B(_04945_),
    .C(_04946_),
    .D(_04943_),
    .Y(_04960_)
  );
  INVX1 _11001_ (
    .A(_04960_),
    .Y(_04961_)
  );
  XNOR2X1 _11002_ (
    .A(_04959_),
    .B(_04961_),
    .Y(_04962_)
  );
  INVX1 _11003_ (
    .A(_04962_),
    .Y(_04963_)
  );
  NAND2X1 _11004_ (
    .A(_04958_),
    .B(_04963_),
    .Y(_04964_)
  );
  XOR2X1 _11005_ (
    .A(_04958_),
    .B(_04962_),
    .Y(_04965_)
  );
  XNOR2X1 _11006_ (
    .A(_04949_),
    .B(_04950_),
    .Y(_04966_)
  );
  OAI21X1 _11007_ (
    .A(_04965_),
    .B(_04966_),
    .C(_04951_),
    .Y(_04967_)
  );
  XOR2X1 _11008_ (
    .A(_04920_),
    .B(_04921_),
    .Y(_04968_)
  );
  NAND2X1 _11009_ (
    .A(_04967_),
    .B(_04968_),
    .Y(_04969_)
  );
  OAI21X1 _11010_ (
    .A(_04959_),
    .B(_04961_),
    .C(_04964_),
    .Y(_04970_)
  );
  INVX1 _11011_ (
    .A(_04970_),
    .Y(_04971_)
  );
  XNOR2X1 _11012_ (
    .A(_04967_),
    .B(_04968_),
    .Y(_04972_)
  );
  OAI21X1 _11013_ (
    .A(_04971_),
    .B(_04972_),
    .C(_04969_),
    .Y(_04973_)
  );
  NAND2X1 _11014_ (
    .A(_04934_),
    .B(_04973_),
    .Y(_04974_)
  );
  NOR2X1 _11015_ (
    .A(_04933_),
    .B(_04974_),
    .Y(_04975_)
  );
  XOR2X1 _11016_ (
    .A(_04933_),
    .B(_04974_),
    .Y(_04976_)
  );
  NAND2X1 _11017_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04638_),
    .Y(_04977_)
  );
  NAND2X1 _11018_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04642_),
    .Y(_04978_)
  );
  NAND2X1 _11019_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04651_),
    .Y(_04979_)
  );
  XNOR2X1 _11020_ (
    .A(_04936_),
    .B(_04977_),
    .Y(_04980_)
  );
  OAI22X1 _11021_ (
    .A(_04935_),
    .B(_04978_),
    .C(_04979_),
    .D(_04980_),
    .Y(_04981_)
  );
  XNOR2X1 _11022_ (
    .A(_04937_),
    .B(_04938_),
    .Y(_04982_)
  );
  INVX1 _11023_ (
    .A(_04982_),
    .Y(_04983_)
  );
  NAND2X1 _11024_ (
    .A(_04981_),
    .B(_04983_),
    .Y(_04984_)
  );
  NAND2X1 _11025_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04657_),
    .Y(_04985_)
  );
  NAND2X1 _11026_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04660_),
    .Y(_04986_)
  );
  NAND2X1 _11027_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04663_),
    .Y(_04987_)
  );
  XNOR2X1 _11028_ (
    .A(_04945_),
    .B(_04986_),
    .Y(_04988_)
  );
  XNOR2X1 _11029_ (
    .A(_04985_),
    .B(_04988_),
    .Y(_04989_)
  );
  XOR2X1 _11030_ (
    .A(_04981_),
    .B(_04982_),
    .Y(_04990_)
  );
  OAI21X1 _11031_ (
    .A(_04989_),
    .B(_04990_),
    .C(_04984_),
    .Y(_04991_)
  );
  XOR2X1 _11032_ (
    .A(_04947_),
    .B(_04948_),
    .Y(_04992_)
  );
  NAND2X1 _11033_ (
    .A(_04991_),
    .B(_04992_),
    .Y(_04993_)
  );
  NAND2X1 _11034_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04685_),
    .Y(_04994_)
  );
  NAND2X1 _11035_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04688_),
    .Y(_04995_)
  );
  NOR2X1 _11036_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04693_),
    .Y(_04996_)
  );
  INVX1 _11037_ (
    .A(_04996_),
    .Y(_04997_)
  );
  NAND2X1 _11038_ (
    .A(_04953_),
    .B(_04994_),
    .Y(_04998_)
  );
  OAI21X1 _11039_ (
    .A(_04952_),
    .B(_04995_),
    .C(_04998_),
    .Y(_04999_)
  );
  OAI22X1 _11040_ (
    .A(_04952_),
    .B(_04995_),
    .C(_04997_),
    .D(_04999_),
    .Y(_05000_)
  );
  XNOR2X1 _11041_ (
    .A(_04955_),
    .B(_04957_),
    .Y(_05001_)
  );
  OAI22X1 _11042_ (
    .A(_04944_),
    .B(_04987_),
    .C(_04988_),
    .D(_04985_),
    .Y(_05002_)
  );
  INVX1 _11043_ (
    .A(_05002_),
    .Y(_05003_)
  );
  XNOR2X1 _11044_ (
    .A(_05001_),
    .B(_05003_),
    .Y(_05004_)
  );
  INVX1 _11045_ (
    .A(_05004_),
    .Y(_05005_)
  );
  NAND2X1 _11046_ (
    .A(_05000_),
    .B(_05005_),
    .Y(_05006_)
  );
  XOR2X1 _11047_ (
    .A(_05000_),
    .B(_05004_),
    .Y(_05007_)
  );
  XNOR2X1 _11048_ (
    .A(_04991_),
    .B(_04992_),
    .Y(_05008_)
  );
  OAI21X1 _11049_ (
    .A(_05007_),
    .B(_05008_),
    .C(_04993_),
    .Y(_05009_)
  );
  XOR2X1 _11050_ (
    .A(_04965_),
    .B(_04966_),
    .Y(_05010_)
  );
  NAND2X1 _11051_ (
    .A(_05009_),
    .B(_05010_),
    .Y(_05011_)
  );
  OAI21X1 _11052_ (
    .A(_05001_),
    .B(_05003_),
    .C(_05006_),
    .Y(_05012_)
  );
  INVX1 _11053_ (
    .A(_05012_),
    .Y(_05013_)
  );
  XNOR2X1 _11054_ (
    .A(_05009_),
    .B(_05010_),
    .Y(_05014_)
  );
  OAI21X1 _11055_ (
    .A(_05013_),
    .B(_05014_),
    .C(_05011_),
    .Y(_05015_)
  );
  XNOR2X1 _11056_ (
    .A(_04970_),
    .B(_04972_),
    .Y(_05016_)
  );
  NAND2X1 _11057_ (
    .A(_05015_),
    .B(_05016_),
    .Y(_05017_)
  );
  XNOR2X1 _11058_ (
    .A(_04934_),
    .B(_04973_),
    .Y(_05018_)
  );
  OR2X1 _11059_ (
    .A(_05017_),
    .B(_05018_),
    .Y(_05019_)
  );
  XOR2X1 _11060_ (
    .A(_05017_),
    .B(_05018_),
    .Y(_05020_)
  );
  INVX1 _11061_ (
    .A(_05020_),
    .Y(_05021_)
  );
  NAND2X1 _11062_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04638_),
    .Y(_05022_)
  );
  NAND2X1 _11063_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04642_),
    .Y(_05023_)
  );
  NAND2X1 _11064_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04651_),
    .Y(_05024_)
  );
  XNOR2X1 _11065_ (
    .A(_04978_),
    .B(_05022_),
    .Y(_05025_)
  );
  OAI22X1 _11066_ (
    .A(_04977_),
    .B(_05023_),
    .C(_05024_),
    .D(_05025_),
    .Y(_05026_)
  );
  XNOR2X1 _11067_ (
    .A(_04979_),
    .B(_04980_),
    .Y(_05027_)
  );
  INVX1 _11068_ (
    .A(_05027_),
    .Y(_05028_)
  );
  NAND2X1 _11069_ (
    .A(_05026_),
    .B(_05028_),
    .Y(_05029_)
  );
  NAND2X1 _11070_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04657_),
    .Y(_05030_)
  );
  NAND2X1 _11071_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04660_),
    .Y(_05031_)
  );
  NAND2X1 _11072_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04663_),
    .Y(_05032_)
  );
  XNOR2X1 _11073_ (
    .A(_04987_),
    .B(_05031_),
    .Y(_05033_)
  );
  XNOR2X1 _11074_ (
    .A(_05030_),
    .B(_05033_),
    .Y(_05034_)
  );
  XOR2X1 _11075_ (
    .A(_05026_),
    .B(_05027_),
    .Y(_05035_)
  );
  OAI21X1 _11076_ (
    .A(_05034_),
    .B(_05035_),
    .C(_05029_),
    .Y(_05036_)
  );
  XOR2X1 _11077_ (
    .A(_04989_),
    .B(_04990_),
    .Y(_05037_)
  );
  NAND2X1 _11078_ (
    .A(_05036_),
    .B(_05037_),
    .Y(_05038_)
  );
  NAND2X1 _11079_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04685_),
    .Y(_05039_)
  );
  NAND2X1 _11080_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04688_),
    .Y(_05040_)
  );
  NOR2X1 _11081_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04693_),
    .Y(_05041_)
  );
  INVX1 _11082_ (
    .A(_05041_),
    .Y(_05042_)
  );
  NAND2X1 _11083_ (
    .A(_04995_),
    .B(_05039_),
    .Y(_05043_)
  );
  OAI21X1 _11084_ (
    .A(_04994_),
    .B(_05040_),
    .C(_05043_),
    .Y(_05044_)
  );
  OAI22X1 _11085_ (
    .A(_04994_),
    .B(_05040_),
    .C(_05042_),
    .D(_05044_),
    .Y(_05045_)
  );
  XNOR2X1 _11086_ (
    .A(_04997_),
    .B(_04999_),
    .Y(_05046_)
  );
  OAI22X1 _11087_ (
    .A(_04986_),
    .B(_05032_),
    .C(_05033_),
    .D(_05030_),
    .Y(_05047_)
  );
  INVX1 _11088_ (
    .A(_05047_),
    .Y(_05048_)
  );
  XNOR2X1 _11089_ (
    .A(_05046_),
    .B(_05048_),
    .Y(_05049_)
  );
  INVX1 _11090_ (
    .A(_05049_),
    .Y(_05050_)
  );
  NAND2X1 _11091_ (
    .A(_05045_),
    .B(_05050_),
    .Y(_05051_)
  );
  XOR2X1 _11092_ (
    .A(_05045_),
    .B(_05049_),
    .Y(_05052_)
  );
  XNOR2X1 _11093_ (
    .A(_05036_),
    .B(_05037_),
    .Y(_05053_)
  );
  OAI21X1 _11094_ (
    .A(_05052_),
    .B(_05053_),
    .C(_05038_),
    .Y(_05054_)
  );
  XOR2X1 _11095_ (
    .A(_05007_),
    .B(_05008_),
    .Y(_05055_)
  );
  NAND2X1 _11096_ (
    .A(_05054_),
    .B(_05055_),
    .Y(_05056_)
  );
  OAI21X1 _11097_ (
    .A(_05046_),
    .B(_05048_),
    .C(_05051_),
    .Y(_05057_)
  );
  INVX1 _11098_ (
    .A(_05057_),
    .Y(_05058_)
  );
  XNOR2X1 _11099_ (
    .A(_05054_),
    .B(_05055_),
    .Y(_05059_)
  );
  OAI21X1 _11100_ (
    .A(_05058_),
    .B(_05059_),
    .C(_05056_),
    .Y(_05060_)
  );
  XNOR2X1 _11101_ (
    .A(_05012_),
    .B(_05014_),
    .Y(_05061_)
  );
  NAND2X1 _11102_ (
    .A(_05060_),
    .B(_05061_),
    .Y(_05062_)
  );
  XNOR2X1 _11103_ (
    .A(_05015_),
    .B(_05016_),
    .Y(_05063_)
  );
  NOR2X1 _11104_ (
    .A(_05062_),
    .B(_05063_),
    .Y(_05064_)
  );
  NAND2X1 _11105_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04638_),
    .Y(_05065_)
  );
  NAND2X1 _11106_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04642_),
    .Y(_05066_)
  );
  NAND2X1 _11107_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04651_),
    .Y(_05067_)
  );
  XNOR2X1 _11108_ (
    .A(_05023_),
    .B(_05065_),
    .Y(_05068_)
  );
  OAI22X1 _11109_ (
    .A(_05022_),
    .B(_05066_),
    .C(_05067_),
    .D(_05068_),
    .Y(_05069_)
  );
  XNOR2X1 _11110_ (
    .A(_05024_),
    .B(_05025_),
    .Y(_05070_)
  );
  INVX1 _11111_ (
    .A(_05070_),
    .Y(_05071_)
  );
  NAND2X1 _11112_ (
    .A(_05069_),
    .B(_05071_),
    .Y(_05072_)
  );
  NAND2X1 _11113_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04657_),
    .Y(_05073_)
  );
  NAND2X1 _11114_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04660_),
    .Y(_05074_)
  );
  NAND2X1 _11115_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04663_),
    .Y(_05075_)
  );
  XNOR2X1 _11116_ (
    .A(_05032_),
    .B(_05074_),
    .Y(_05076_)
  );
  XNOR2X1 _11117_ (
    .A(_05073_),
    .B(_05076_),
    .Y(_05077_)
  );
  XOR2X1 _11118_ (
    .A(_05069_),
    .B(_05070_),
    .Y(_05078_)
  );
  OAI21X1 _11119_ (
    .A(_05077_),
    .B(_05078_),
    .C(_05072_),
    .Y(_05079_)
  );
  XOR2X1 _11120_ (
    .A(_05034_),
    .B(_05035_),
    .Y(_05080_)
  );
  NAND2X1 _11121_ (
    .A(_05079_),
    .B(_05080_),
    .Y(_05081_)
  );
  NAND2X1 _11122_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04685_),
    .Y(_05082_)
  );
  NAND2X1 _11123_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04688_),
    .Y(_05083_)
  );
  NOR2X1 _11124_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04693_),
    .Y(_05084_)
  );
  INVX1 _11125_ (
    .A(_05084_),
    .Y(_05085_)
  );
  NAND2X1 _11126_ (
    .A(_05040_),
    .B(_05082_),
    .Y(_05086_)
  );
  OAI21X1 _11127_ (
    .A(_05039_),
    .B(_05083_),
    .C(_05086_),
    .Y(_05087_)
  );
  OAI22X1 _11128_ (
    .A(_05039_),
    .B(_05083_),
    .C(_05085_),
    .D(_05087_),
    .Y(_05088_)
  );
  XNOR2X1 _11129_ (
    .A(_05042_),
    .B(_05044_),
    .Y(_05089_)
  );
  OAI22X1 _11130_ (
    .A(_05031_),
    .B(_05075_),
    .C(_05076_),
    .D(_05073_),
    .Y(_05090_)
  );
  INVX1 _11131_ (
    .A(_05090_),
    .Y(_05091_)
  );
  XNOR2X1 _11132_ (
    .A(_05089_),
    .B(_05091_),
    .Y(_05092_)
  );
  INVX1 _11133_ (
    .A(_05092_),
    .Y(_05093_)
  );
  NAND2X1 _11134_ (
    .A(_05088_),
    .B(_05093_),
    .Y(_05094_)
  );
  XOR2X1 _11135_ (
    .A(_05088_),
    .B(_05092_),
    .Y(_05095_)
  );
  XNOR2X1 _11136_ (
    .A(_05079_),
    .B(_05080_),
    .Y(_05096_)
  );
  OAI21X1 _11137_ (
    .A(_05095_),
    .B(_05096_),
    .C(_05081_),
    .Y(_05097_)
  );
  XOR2X1 _11138_ (
    .A(_05052_),
    .B(_05053_),
    .Y(_05098_)
  );
  NAND2X1 _11139_ (
    .A(_05097_),
    .B(_05098_),
    .Y(_05099_)
  );
  OAI21X1 _11140_ (
    .A(_05089_),
    .B(_05091_),
    .C(_05094_),
    .Y(_05100_)
  );
  INVX1 _11141_ (
    .A(_05100_),
    .Y(_05101_)
  );
  XNOR2X1 _11142_ (
    .A(_05097_),
    .B(_05098_),
    .Y(_05102_)
  );
  OAI21X1 _11143_ (
    .A(_05101_),
    .B(_05102_),
    .C(_05099_),
    .Y(_05103_)
  );
  XNOR2X1 _11144_ (
    .A(_05057_),
    .B(_05059_),
    .Y(_05104_)
  );
  NAND2X1 _11145_ (
    .A(_05103_),
    .B(_05104_),
    .Y(_05105_)
  );
  XNOR2X1 _11146_ (
    .A(_05060_),
    .B(_05061_),
    .Y(_05106_)
  );
  NOR2X1 _11147_ (
    .A(_05105_),
    .B(_05106_),
    .Y(_05107_)
  );
  OR2X1 _11148_ (
    .A(_05105_),
    .B(_05106_),
    .Y(_05108_)
  );
  AND2X1 _11149_ (
    .A(_05105_),
    .B(_05106_),
    .Y(_05109_)
  );
  NOR2X1 _11150_ (
    .A(_05107_),
    .B(_05109_),
    .Y(_05110_)
  );
  OR2X1 _11151_ (
    .A(_04611_),
    .B(_04641_),
    .Y(_05111_)
  );
  NOR2X1 _11152_ (
    .A(_05065_),
    .B(_05111_),
    .Y(_05112_)
  );
  NAND2X1 _11153_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04651_),
    .Y(_05113_)
  );
  OAI21X1 _11154_ (
    .A(_04611_),
    .B(_04637_),
    .C(_05066_),
    .Y(_05114_)
  );
  OAI21X1 _11155_ (
    .A(_05065_),
    .B(_05111_),
    .C(_05114_),
    .Y(_05115_)
  );
  NOR2X1 _11156_ (
    .A(_05113_),
    .B(_05115_),
    .Y(_05116_)
  );
  NOR2X1 _11157_ (
    .A(_05112_),
    .B(_05116_),
    .Y(_05117_)
  );
  XNOR2X1 _11158_ (
    .A(_05067_),
    .B(_05068_),
    .Y(_05118_)
  );
  NOR2X1 _11159_ (
    .A(_05117_),
    .B(_05118_),
    .Y(_05119_)
  );
  NAND2X1 _11160_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04657_),
    .Y(_05120_)
  );
  NAND2X1 _11161_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04660_),
    .Y(_05121_)
  );
  AND2X1 _11162_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04663_),
    .Y(_05122_)
  );
  OR2X1 _11163_ (
    .A(_05075_),
    .B(_05121_),
    .Y(_05123_)
  );
  XNOR2X1 _11164_ (
    .A(_05075_),
    .B(_05121_),
    .Y(_05124_)
  );
  XNOR2X1 _11165_ (
    .A(_05120_),
    .B(_05124_),
    .Y(_05125_)
  );
  INVX1 _11166_ (
    .A(_05125_),
    .Y(_05126_)
  );
  XOR2X1 _11167_ (
    .A(_05117_),
    .B(_05118_),
    .Y(_05127_)
  );
  AOI21X1 _11168_ (
    .A(_05126_),
    .B(_05127_),
    .C(_05119_),
    .Y(_05128_)
  );
  INVX1 _11169_ (
    .A(_05128_),
    .Y(_05129_)
  );
  XOR2X1 _11170_ (
    .A(_05077_),
    .B(_05078_),
    .Y(_05130_)
  );
  NAND2X1 _11171_ (
    .A(_05129_),
    .B(_05130_),
    .Y(_05131_)
  );
  NAND2X1 _11172_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04685_),
    .Y(_05132_)
  );
  NAND2X1 _11173_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04688_),
    .Y(_05133_)
  );
  NOR2X1 _11174_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04693_),
    .Y(_05134_)
  );
  INVX1 _11175_ (
    .A(_05134_),
    .Y(_05135_)
  );
  NAND2X1 _11176_ (
    .A(_05083_),
    .B(_05132_),
    .Y(_05136_)
  );
  OAI21X1 _11177_ (
    .A(_05082_),
    .B(_05133_),
    .C(_05136_),
    .Y(_05137_)
  );
  OAI22X1 _11178_ (
    .A(_05082_),
    .B(_05133_),
    .C(_05135_),
    .D(_05137_),
    .Y(_05138_)
  );
  XNOR2X1 _11179_ (
    .A(_05085_),
    .B(_05087_),
    .Y(_05139_)
  );
  INVX1 _11180_ (
    .A(_05139_),
    .Y(_05140_)
  );
  OAI21X1 _11181_ (
    .A(_05120_),
    .B(_05124_),
    .C(_05123_),
    .Y(_05141_)
  );
  AND2X1 _11182_ (
    .A(_05140_),
    .B(_05141_),
    .Y(_05142_)
  );
  XOR2X1 _11183_ (
    .A(_05139_),
    .B(_05141_),
    .Y(_05143_)
  );
  INVX1 _11184_ (
    .A(_05143_),
    .Y(_05144_)
  );
  XOR2X1 _11185_ (
    .A(_05138_),
    .B(_05143_),
    .Y(_05145_)
  );
  NOR2X1 _11186_ (
    .A(_05129_),
    .B(_05130_),
    .Y(_05146_)
  );
  XNOR2X1 _11187_ (
    .A(_05128_),
    .B(_05130_),
    .Y(_05147_)
  );
  OAI21X1 _11188_ (
    .A(_05145_),
    .B(_05146_),
    .C(_05131_),
    .Y(_05148_)
  );
  XOR2X1 _11189_ (
    .A(_05095_),
    .B(_05096_),
    .Y(_05149_)
  );
  NAND2X1 _11190_ (
    .A(_05148_),
    .B(_05149_),
    .Y(_05150_)
  );
  AOI21X1 _11191_ (
    .A(_05138_),
    .B(_05144_),
    .C(_05142_),
    .Y(_05151_)
  );
  XNOR2X1 _11192_ (
    .A(_05148_),
    .B(_05149_),
    .Y(_05152_)
  );
  OAI21X1 _11193_ (
    .A(_05151_),
    .B(_05152_),
    .C(_05150_),
    .Y(_05153_)
  );
  XNOR2X1 _11194_ (
    .A(_05100_),
    .B(_05102_),
    .Y(_05154_)
  );
  NAND2X1 _11195_ (
    .A(_05153_),
    .B(_05154_),
    .Y(_05155_)
  );
  XNOR2X1 _11196_ (
    .A(_05103_),
    .B(_05104_),
    .Y(_05156_)
  );
  NOR2X1 _11197_ (
    .A(_05155_),
    .B(_05156_),
    .Y(_05157_)
  );
  XOR2X1 _11198_ (
    .A(_05155_),
    .B(_05156_),
    .Y(_05158_)
  );
  NOR2X1 _11199_ (
    .A(_04609_),
    .B(_04637_),
    .Y(_05159_)
  );
  XOR2X1 _11200_ (
    .A(_04693_),
    .B(_05111_),
    .Y(_05160_)
  );
  NAND2X1 _11201_ (
    .A(_05159_),
    .B(_05160_),
    .Y(_05161_)
  );
  OAI21X1 _11202_ (
    .A(_04693_),
    .B(_05111_),
    .C(_05161_),
    .Y(_05162_)
  );
  XNOR2X1 _11203_ (
    .A(_05113_),
    .B(_05115_),
    .Y(_05163_)
  );
  INVX1 _11204_ (
    .A(_05163_),
    .Y(_05164_)
  );
  NAND2X1 _11205_ (
    .A(_05162_),
    .B(_05164_),
    .Y(_05165_)
  );
  NAND2X1 _11206_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04657_),
    .Y(_05166_)
  );
  NAND2X1 _11207_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04660_),
    .Y(_05167_)
  );
  NAND2X1 _11208_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04663_),
    .Y(_05168_)
  );
  XOR2X1 _11209_ (
    .A(_05122_),
    .B(_05167_),
    .Y(_05169_)
  );
  XNOR2X1 _11210_ (
    .A(_05166_),
    .B(_05169_),
    .Y(_05170_)
  );
  XOR2X1 _11211_ (
    .A(_05162_),
    .B(_05163_),
    .Y(_05171_)
  );
  OAI21X1 _11212_ (
    .A(_05170_),
    .B(_05171_),
    .C(_05165_),
    .Y(_05172_)
  );
  XNOR2X1 _11213_ (
    .A(_05125_),
    .B(_05127_),
    .Y(_05173_)
  );
  NAND2X1 _11214_ (
    .A(_05172_),
    .B(_05173_),
    .Y(_05174_)
  );
  NAND2X1 _11215_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04685_),
    .Y(_05175_)
  );
  NAND2X1 _11216_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04688_),
    .Y(_05176_)
  );
  OR2X1 _11217_ (
    .A(_05132_),
    .B(_05176_),
    .Y(_05177_)
  );
  NOR2X1 _11218_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04693_),
    .Y(_05178_)
  );
  NAND2X1 _11219_ (
    .A(_05133_),
    .B(_05175_),
    .Y(_05179_)
  );
  OAI21X1 _11220_ (
    .A(_05132_),
    .B(_05176_),
    .C(_05179_),
    .Y(_05180_)
  );
  NAND3X1 _11221_ (
    .A(_05177_),
    .B(_05178_),
    .C(_05179_),
    .Y(_05181_)
  );
  OAI21X1 _11222_ (
    .A(_05132_),
    .B(_05176_),
    .C(_05181_),
    .Y(_05182_)
  );
  XNOR2X1 _11223_ (
    .A(_05135_),
    .B(_05137_),
    .Y(_05183_)
  );
  INVX1 _11224_ (
    .A(_05183_),
    .Y(_05184_)
  );
  OAI22X1 _11225_ (
    .A(_05121_),
    .B(_05168_),
    .C(_05169_),
    .D(_05166_),
    .Y(_05185_)
  );
  XOR2X1 _11226_ (
    .A(_05183_),
    .B(_05185_),
    .Y(_05186_)
  );
  AOI21X1 _11227_ (
    .A(_05177_),
    .B(_05181_),
    .C(_05186_),
    .Y(_05187_)
  );
  XOR2X1 _11228_ (
    .A(_05182_),
    .B(_05186_),
    .Y(_05188_)
  );
  XNOR2X1 _11229_ (
    .A(_05172_),
    .B(_05173_),
    .Y(_05189_)
  );
  OAI21X1 _11230_ (
    .A(_05188_),
    .B(_05189_),
    .C(_05174_),
    .Y(_05190_)
  );
  XNOR2X1 _11231_ (
    .A(_05145_),
    .B(_05147_),
    .Y(_05191_)
  );
  NAND2X1 _11232_ (
    .A(_05190_),
    .B(_05191_),
    .Y(_05192_)
  );
  AOI21X1 _11233_ (
    .A(_05184_),
    .B(_05185_),
    .C(_05187_),
    .Y(_05193_)
  );
  XNOR2X1 _11234_ (
    .A(_05190_),
    .B(_05191_),
    .Y(_05194_)
  );
  OAI21X1 _11235_ (
    .A(_05193_),
    .B(_05194_),
    .C(_05192_),
    .Y(_05195_)
  );
  XOR2X1 _11236_ (
    .A(_05151_),
    .B(_05152_),
    .Y(_05196_)
  );
  NAND2X1 _11237_ (
    .A(_05195_),
    .B(_05196_),
    .Y(_05197_)
  );
  XNOR2X1 _11238_ (
    .A(_05153_),
    .B(_05154_),
    .Y(_05198_)
  );
  OR2X1 _11239_ (
    .A(_05197_),
    .B(_05198_),
    .Y(_05199_)
  );
  XOR2X1 _11240_ (
    .A(_05197_),
    .B(_05198_),
    .Y(_05200_)
  );
  INVX1 _11241_ (
    .A(_05200_),
    .Y(_05201_)
  );
  NOR2X1 _11242_ (
    .A(_04607_),
    .B(_04637_),
    .Y(_05202_)
  );
  NOR2X1 _11243_ (
    .A(_04609_),
    .B(_04641_),
    .Y(_05203_)
  );
  NOR2X1 _11244_ (
    .A(_04607_),
    .B(_04641_),
    .Y(_05204_)
  );
  AND2X1 _11245_ (
    .A(_05159_),
    .B(_05204_),
    .Y(_05205_)
  );
  AND2X1 _11246_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04651_),
    .Y(_05206_)
  );
  OR2X1 _11247_ (
    .A(_05202_),
    .B(_05203_),
    .Y(_05207_)
  );
  XNOR2X1 _11248_ (
    .A(_05202_),
    .B(_05203_),
    .Y(_05208_)
  );
  AOI21X1 _11249_ (
    .A(_05206_),
    .B(_05207_),
    .C(_05205_),
    .Y(_05209_)
  );
  XNOR2X1 _11250_ (
    .A(_05159_),
    .B(_05160_),
    .Y(_05210_)
  );
  NAND2X1 _11251_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04660_),
    .Y(_05211_)
  );
  NAND2X1 _11252_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04651_),
    .Y(_05212_)
  );
  NAND2X1 _11253_ (
    .A(_05122_),
    .B(_05206_),
    .Y(_05213_)
  );
  XNOR2X1 _11254_ (
    .A(_05168_),
    .B(_05212_),
    .Y(_05214_)
  );
  XNOR2X1 _11255_ (
    .A(_05211_),
    .B(_05214_),
    .Y(_05215_)
  );
  INVX1 _11256_ (
    .A(_05215_),
    .Y(_05216_)
  );
  XOR2X1 _11257_ (
    .A(_05209_),
    .B(_05210_),
    .Y(_05217_)
  );
  NAND2X1 _11258_ (
    .A(_05216_),
    .B(_05217_),
    .Y(_05218_)
  );
  OAI21X1 _11259_ (
    .A(_05209_),
    .B(_05210_),
    .C(_05218_),
    .Y(_05219_)
  );
  XOR2X1 _11260_ (
    .A(_05170_),
    .B(_05171_),
    .Y(_05220_)
  );
  NAND2X1 _11261_ (
    .A(_05219_),
    .B(_05220_),
    .Y(_05221_)
  );
  NAND2X1 _11262_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04657_),
    .Y(_05222_)
  );
  NAND2X1 _11263_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04657_),
    .Y(_05223_)
  );
  NAND2X1 _11264_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04685_),
    .Y(_05224_)
  );
  XNOR2X1 _11265_ (
    .A(_05176_),
    .B(_05222_),
    .Y(_05225_)
  );
  OAI22X1 _11266_ (
    .A(_05133_),
    .B(_05223_),
    .C(_05224_),
    .D(_05225_),
    .Y(_05226_)
  );
  XOR2X1 _11267_ (
    .A(_05178_),
    .B(_05180_),
    .Y(_05227_)
  );
  INVX1 _11268_ (
    .A(_05227_),
    .Y(_05228_)
  );
  OAI21X1 _11269_ (
    .A(_05211_),
    .B(_05214_),
    .C(_05213_),
    .Y(_05229_)
  );
  AND2X1 _11270_ (
    .A(_05228_),
    .B(_05229_),
    .Y(_05230_)
  );
  XOR2X1 _11271_ (
    .A(_05227_),
    .B(_05229_),
    .Y(_05231_)
  );
  INVX1 _11272_ (
    .A(_05231_),
    .Y(_05232_)
  );
  XOR2X1 _11273_ (
    .A(_05226_),
    .B(_05231_),
    .Y(_05233_)
  );
  XNOR2X1 _11274_ (
    .A(_05219_),
    .B(_05220_),
    .Y(_05234_)
  );
  OAI21X1 _11275_ (
    .A(_05233_),
    .B(_05234_),
    .C(_05221_),
    .Y(_05235_)
  );
  XOR2X1 _11276_ (
    .A(_05188_),
    .B(_05189_),
    .Y(_05236_)
  );
  NAND2X1 _11277_ (
    .A(_05235_),
    .B(_05236_),
    .Y(_05237_)
  );
  AOI21X1 _11278_ (
    .A(_05226_),
    .B(_05232_),
    .C(_05230_),
    .Y(_05238_)
  );
  XNOR2X1 _11279_ (
    .A(_05235_),
    .B(_05236_),
    .Y(_05239_)
  );
  OAI21X1 _11280_ (
    .A(_05238_),
    .B(_05239_),
    .C(_05237_),
    .Y(_05240_)
  );
  XOR2X1 _11281_ (
    .A(_05193_),
    .B(_05194_),
    .Y(_05241_)
  );
  NAND2X1 _11282_ (
    .A(_05240_),
    .B(_05241_),
    .Y(_05242_)
  );
  XNOR2X1 _11283_ (
    .A(_05195_),
    .B(_05196_),
    .Y(_05243_)
  );
  NOR2X1 _11284_ (
    .A(_05242_),
    .B(_05243_),
    .Y(_05244_)
  );
  NOR2X1 _11285_ (
    .A(_04605_),
    .B(_04637_),
    .Y(_05245_)
  );
  NOR2X1 _11286_ (
    .A(_04605_),
    .B(_04641_),
    .Y(_05246_)
  );
  NAND2X1 _11287_ (
    .A(_05204_),
    .B(_05245_),
    .Y(_05247_)
  );
  NAND2X1 _11288_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04651_),
    .Y(_05248_)
  );
  NOR2X1 _11289_ (
    .A(_05204_),
    .B(_05245_),
    .Y(_05249_)
  );
  XOR2X1 _11290_ (
    .A(_05204_),
    .B(_05245_),
    .Y(_05250_)
  );
  OAI21X1 _11291_ (
    .A(_05248_),
    .B(_05249_),
    .C(_05247_),
    .Y(_05251_)
  );
  XNOR2X1 _11292_ (
    .A(_05206_),
    .B(_05208_),
    .Y(_05252_)
  );
  NAND2X1 _11293_ (
    .A(_05251_),
    .B(_05252_),
    .Y(_05253_)
  );
  NAND2X1 _11294_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04660_),
    .Y(_05254_)
  );
  NAND2X1 _11295_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04663_),
    .Y(_05255_)
  );
  NAND2X1 _11296_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04663_),
    .Y(_05256_)
  );
  XNOR2X1 _11297_ (
    .A(_05254_),
    .B(_05255_),
    .Y(_05257_)
  );
  XNOR2X1 _11298_ (
    .A(_05223_),
    .B(_05257_),
    .Y(_05258_)
  );
  XNOR2X1 _11299_ (
    .A(_05251_),
    .B(_05252_),
    .Y(_05259_)
  );
  OAI21X1 _11300_ (
    .A(_05258_),
    .B(_05259_),
    .C(_05253_),
    .Y(_05260_)
  );
  XNOR2X1 _11301_ (
    .A(_05215_),
    .B(_05217_),
    .Y(_05261_)
  );
  NAND2X1 _11302_ (
    .A(_05260_),
    .B(_05261_),
    .Y(_05262_)
  );
  AND2X1 _11303_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04688_),
    .Y(_05263_)
  );
  NAND3X1 _11304_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04685_),
    .C(_05263_),
    .Y(_05264_)
  );
  INVX1 _11305_ (
    .A(_05264_),
    .Y(_05265_)
  );
  XNOR2X1 _11306_ (
    .A(_05224_),
    .B(_05225_),
    .Y(_05266_)
  );
  INVX1 _11307_ (
    .A(_05266_),
    .Y(_05267_)
  );
  OAI22X1 _11308_ (
    .A(_05211_),
    .B(_05256_),
    .C(_05257_),
    .D(_05223_),
    .Y(_05268_)
  );
  XOR2X1 _11309_ (
    .A(_05266_),
    .B(_05268_),
    .Y(_05269_)
  );
  NOR2X1 _11310_ (
    .A(_05264_),
    .B(_05269_),
    .Y(_05270_)
  );
  XNOR2X1 _11311_ (
    .A(_05264_),
    .B(_05269_),
    .Y(_05271_)
  );
  XNOR2X1 _11312_ (
    .A(_05260_),
    .B(_05261_),
    .Y(_05272_)
  );
  OAI21X1 _11313_ (
    .A(_05271_),
    .B(_05272_),
    .C(_05262_),
    .Y(_05273_)
  );
  XOR2X1 _11314_ (
    .A(_05233_),
    .B(_05234_),
    .Y(_05274_)
  );
  NAND2X1 _11315_ (
    .A(_05273_),
    .B(_05274_),
    .Y(_05275_)
  );
  AOI21X1 _11316_ (
    .A(_05267_),
    .B(_05268_),
    .C(_05270_),
    .Y(_05276_)
  );
  XNOR2X1 _11317_ (
    .A(_05273_),
    .B(_05274_),
    .Y(_05277_)
  );
  OAI21X1 _11318_ (
    .A(_05276_),
    .B(_05277_),
    .C(_05275_),
    .Y(_05278_)
  );
  XOR2X1 _11319_ (
    .A(_05238_),
    .B(_05239_),
    .Y(_05279_)
  );
  NAND2X1 _11320_ (
    .A(_05278_),
    .B(_05279_),
    .Y(_05280_)
  );
  XNOR2X1 _11321_ (
    .A(_05240_),
    .B(_05241_),
    .Y(_05281_)
  );
  OR2X1 _11322_ (
    .A(_05280_),
    .B(_05281_),
    .Y(_05282_)
  );
  XOR2X1 _11323_ (
    .A(_05280_),
    .B(_05281_),
    .Y(_05283_)
  );
  INVX1 _11324_ (
    .A(_05283_),
    .Y(_05284_)
  );
  NOR2X1 _11325_ (
    .A(_04603_),
    .B(_04637_),
    .Y(_05285_)
  );
  NOR2X1 _11326_ (
    .A(_04603_),
    .B(_04641_),
    .Y(_05286_)
  );
  NAND2X1 _11327_ (
    .A(_05246_),
    .B(_05285_),
    .Y(_05287_)
  );
  NAND2X1 _11328_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04651_),
    .Y(_05288_)
  );
  XNOR2X1 _11329_ (
    .A(_05246_),
    .B(_05285_),
    .Y(_05289_)
  );
  OAI21X1 _11330_ (
    .A(_05288_),
    .B(_05289_),
    .C(_05287_),
    .Y(_05290_)
  );
  XNOR2X1 _11331_ (
    .A(_05248_),
    .B(_05250_),
    .Y(_05291_)
  );
  NAND2X1 _11332_ (
    .A(_05290_),
    .B(_05291_),
    .Y(_05292_)
  );
  NAND2X1 _11333_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04657_),
    .Y(_05293_)
  );
  NAND2X1 _11334_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04660_),
    .Y(_05294_)
  );
  AND2X1 _11335_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04663_),
    .Y(_05295_)
  );
  OR2X1 _11336_ (
    .A(_05256_),
    .B(_05294_),
    .Y(_05296_)
  );
  XNOR2X1 _11337_ (
    .A(_05256_),
    .B(_05294_),
    .Y(_05297_)
  );
  XNOR2X1 _11338_ (
    .A(_05293_),
    .B(_05297_),
    .Y(_05298_)
  );
  XNOR2X1 _11339_ (
    .A(_05290_),
    .B(_05291_),
    .Y(_05299_)
  );
  OAI21X1 _11340_ (
    .A(_05298_),
    .B(_05299_),
    .C(_05292_),
    .Y(_05300_)
  );
  XOR2X1 _11341_ (
    .A(_05258_),
    .B(_05259_),
    .Y(_05301_)
  );
  NAND2X1 _11342_ (
    .A(_05300_),
    .B(_05301_),
    .Y(_05302_)
  );
  AOI22X1 _11343_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04685_),
    .C(_04688_),
    .D( multiplier_0.op1_1_ ),
    .Y(_05303_)
  );
  NOR2X1 _11344_ (
    .A(_05265_),
    .B(_05303_),
    .Y(_05304_)
  );
  OAI21X1 _11345_ (
    .A(_05293_),
    .B(_05297_),
    .C(_05296_),
    .Y(_05305_)
  );
  NAND2X1 _11346_ (
    .A(_05304_),
    .B(_05305_),
    .Y(_05306_)
  );
  XNOR2X1 _11347_ (
    .A(_05304_),
    .B(_05305_),
    .Y(_05307_)
  );
  XNOR2X1 _11348_ (
    .A(_05300_),
    .B(_05301_),
    .Y(_05308_)
  );
  OAI21X1 _11349_ (
    .A(_05307_),
    .B(_05308_),
    .C(_05302_),
    .Y(_05309_)
  );
  XNOR2X1 _11350_ (
    .A(_05271_),
    .B(_05272_),
    .Y(_05310_)
  );
  INVX1 _11351_ (
    .A(_05310_),
    .Y(_05311_)
  );
  NAND2X1 _11352_ (
    .A(_05309_),
    .B(_05311_),
    .Y(_05312_)
  );
  XOR2X1 _11353_ (
    .A(_05309_),
    .B(_05310_),
    .Y(_05313_)
  );
  OAI21X1 _11354_ (
    .A(_05306_),
    .B(_05313_),
    .C(_05312_),
    .Y(_05314_)
  );
  XNOR2X1 _11355_ (
    .A(_05276_),
    .B(_05277_),
    .Y(_05315_)
  );
  INVX1 _11356_ (
    .A(_05315_),
    .Y(_05316_)
  );
  NAND2X1 _11357_ (
    .A(_05314_),
    .B(_05316_),
    .Y(_05317_)
  );
  XNOR2X1 _11358_ (
    .A(_05278_),
    .B(_05279_),
    .Y(_05318_)
  );
  NOR2X1 _11359_ (
    .A(_05317_),
    .B(_05318_),
    .Y(_05319_)
  );
  XOR2X1 _11360_ (
    .A(_05317_),
    .B(_05318_),
    .Y(_05320_)
  );
  NOR2X1 _11361_ (
    .A(_04601_),
    .B(_04637_),
    .Y(_05321_)
  );
  NOR2X1 _11362_ (
    .A(_04601_),
    .B(_04641_),
    .Y(_05322_)
  );
  NAND2X1 _11363_ (
    .A(_05286_),
    .B(_05321_),
    .Y(_05323_)
  );
  NAND2X1 _11364_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04651_),
    .Y(_05324_)
  );
  XNOR2X1 _11365_ (
    .A(_05286_),
    .B(_05321_),
    .Y(_05325_)
  );
  OAI21X1 _11366_ (
    .A(_05324_),
    .B(_05325_),
    .C(_05323_),
    .Y(_05326_)
  );
  XOR2X1 _11367_ (
    .A(_05288_),
    .B(_05289_),
    .Y(_05327_)
  );
  NAND2X1 _11368_ (
    .A(_05326_),
    .B(_05327_),
    .Y(_05328_)
  );
  NAND2X1 _11369_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04657_),
    .Y(_05329_)
  );
  NAND2X1 _11370_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04660_),
    .Y(_05330_)
  );
  NAND3X1 _11371_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04660_),
    .C(_05295_),
    .Y(_05331_)
  );
  XOR2X1 _11372_ (
    .A(_05295_),
    .B(_05330_),
    .Y(_05332_)
  );
  XNOR2X1 _11373_ (
    .A(_05329_),
    .B(_05332_),
    .Y(_05333_)
  );
  XNOR2X1 _11374_ (
    .A(_05326_),
    .B(_05327_),
    .Y(_05334_)
  );
  OAI21X1 _11375_ (
    .A(_05333_),
    .B(_05334_),
    .C(_05328_),
    .Y(_05335_)
  );
  XOR2X1 _11376_ (
    .A(_05298_),
    .B(_05299_),
    .Y(_05336_)
  );
  NAND2X1 _11377_ (
    .A(_05335_),
    .B(_05336_),
    .Y(_05337_)
  );
  OAI21X1 _11378_ (
    .A(_05329_),
    .B(_05332_),
    .C(_05331_),
    .Y(_05338_)
  );
  NAND2X1 _11379_ (
    .A(_05263_),
    .B(_05338_),
    .Y(_05339_)
  );
  XNOR2X1 _11380_ (
    .A(_05263_),
    .B(_05338_),
    .Y(_05340_)
  );
  XNOR2X1 _11381_ (
    .A(_05335_),
    .B(_05336_),
    .Y(_05341_)
  );
  OAI21X1 _11382_ (
    .A(_05340_),
    .B(_05341_),
    .C(_05337_),
    .Y(_05342_)
  );
  XOR2X1 _11383_ (
    .A(_05307_),
    .B(_05308_),
    .Y(_05343_)
  );
  NAND2X1 _11384_ (
    .A(_05342_),
    .B(_05343_),
    .Y(_05344_)
  );
  XNOR2X1 _11385_ (
    .A(_05342_),
    .B(_05343_),
    .Y(_05345_)
  );
  OAI21X1 _11386_ (
    .A(_05339_),
    .B(_05345_),
    .C(_05344_),
    .Y(_05346_)
  );
  XOR2X1 _11387_ (
    .A(_05306_),
    .B(_05313_),
    .Y(_05347_)
  );
  NAND2X1 _11388_ (
    .A(_05346_),
    .B(_05347_),
    .Y(_05348_)
  );
  OR2X1 _11389_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04693_),
    .Y(_05349_)
  );
  XNOR2X1 _11390_ (
    .A(_05346_),
    .B(_05347_),
    .Y(_05350_)
  );
  OAI21X1 _11391_ (
    .A(_05349_),
    .B(_05350_),
    .C(_05348_),
    .Y(_05351_)
  );
  XNOR2X1 _11392_ (
    .A(_05314_),
    .B(_05315_),
    .Y(_05352_)
  );
  NAND2X1 _11393_ (
    .A(_05351_),
    .B(_05352_),
    .Y(_05353_)
  );
  XNOR2X1 _11394_ (
    .A(_05351_),
    .B(_05352_),
    .Y(_05354_)
  );
  NAND3X1 _11395_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04638_),
    .C(_05322_),
    .Y(_05355_)
  );
  NAND2X1 _11396_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04651_),
    .Y(_05356_)
  );
  AOI21X1 _11397_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04638_),
    .C(_05322_),
    .Y(_05357_)
  );
  OAI22X1 _11398_ (
    .A(_04599_),
    .B(_04637_),
    .C(_04641_),
    .D(_04601_),
    .Y(_05358_)
  );
  NAND2X1 _11399_ (
    .A(_05355_),
    .B(_05358_),
    .Y(_05359_)
  );
  OAI21X1 _11400_ (
    .A(_05356_),
    .B(_05357_),
    .C(_05355_),
    .Y(_05360_)
  );
  XOR2X1 _11401_ (
    .A(_05324_),
    .B(_05325_),
    .Y(_05361_)
  );
  AND2X1 _11402_ (
    .A(_05360_),
    .B(_05361_),
    .Y(_05362_)
  );
  AOI22X1 _11403_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04660_),
    .C(_04663_),
    .D( multiplier_0.op1_1_ ),
    .Y(_05363_)
  );
  NAND2X1 _11404_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04663_),
    .Y(_05364_)
  );
  NOR2X1 _11405_ (
    .A(_05330_),
    .B(_05364_),
    .Y(_05365_)
  );
  OR2X1 _11406_ (
    .A(_05330_),
    .B(_05364_),
    .Y(_05366_)
  );
  OR2X1 _11407_ (
    .A(_05363_),
    .B(_05365_),
    .Y(_05367_)
  );
  XNOR2X1 _11408_ (
    .A(_05360_),
    .B(_05361_),
    .Y(_05368_)
  );
  NOR2X1 _11409_ (
    .A(_05367_),
    .B(_05368_),
    .Y(_05369_)
  );
  OR2X1 _11410_ (
    .A(_05362_),
    .B(_05369_),
    .Y(_05370_)
  );
  XOR2X1 _11411_ (
    .A(_05333_),
    .B(_05334_),
    .Y(_05371_)
  );
  OAI21X1 _11412_ (
    .A(_05362_),
    .B(_05369_),
    .C(_05371_),
    .Y(_05372_)
  );
  XNOR2X1 _11413_ (
    .A(_05370_),
    .B(_05371_),
    .Y(_05373_)
  );
  OAI21X1 _11414_ (
    .A(_05366_),
    .B(_05373_),
    .C(_05372_),
    .Y(_05374_)
  );
  XOR2X1 _11415_ (
    .A(_05340_),
    .B(_05341_),
    .Y(_05375_)
  );
  NAND2X1 _11416_ (
    .A(_05374_),
    .B(_05375_),
    .Y(_05376_)
  );
  XNOR2X1 _11417_ (
    .A(_05339_),
    .B(_05345_),
    .Y(_05377_)
  );
  OR2X1 _11418_ (
    .A(_05376_),
    .B(_05377_),
    .Y(_05378_)
  );
  XNOR2X1 _11419_ (
    .A(_05349_),
    .B(_05350_),
    .Y(_05379_)
  );
  NOR2X1 _11420_ (
    .A(_05378_),
    .B(_05379_),
    .Y(_05380_)
  );
  NOR2X1 _11421_ (
    .A(_04596_),
    .B(_04637_),
    .Y(_05381_)
  );
  NAND3X1 _11422_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04642_),
    .C(_05381_),
    .Y(_05382_)
  );
  NAND2X1 _11423_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04651_),
    .Y(_05383_)
  );
  OAI22X1 _11424_ (
    .A(_04596_),
    .B(_04637_),
    .C(_04641_),
    .D(_04599_),
    .Y(_05384_)
  );
  NAND2X1 _11425_ (
    .A(_05382_),
    .B(_05384_),
    .Y(_05385_)
  );
  OAI21X1 _11426_ (
    .A(_05383_),
    .B(_05385_),
    .C(_05382_),
    .Y(_05386_)
  );
  XOR2X1 _11427_ (
    .A(_05356_),
    .B(_05359_),
    .Y(_05387_)
  );
  NAND2X1 _11428_ (
    .A(_05386_),
    .B(_05387_),
    .Y(_05388_)
  );
  XNOR2X1 _11429_ (
    .A(_05386_),
    .B(_05387_),
    .Y(_05389_)
  );
  OAI21X1 _11430_ (
    .A(_05364_),
    .B(_05389_),
    .C(_05388_),
    .Y(_05390_)
  );
  XOR2X1 _11431_ (
    .A(_05367_),
    .B(_05368_),
    .Y(_05391_)
  );
  NAND2X1 _11432_ (
    .A(_05390_),
    .B(_05391_),
    .Y(_05392_)
  );
  XNOR2X1 _11433_ (
    .A(_05366_),
    .B(_05373_),
    .Y(_05393_)
  );
  OR2X1 _11434_ (
    .A(_05392_),
    .B(_05393_),
    .Y(_05394_)
  );
  XNOR2X1 _11435_ (
    .A(_05374_),
    .B(_05375_),
    .Y(_04013_)
  );
  NOR2X1 _11436_ (
    .A(_05394_),
    .B(_04013_),
    .Y(_04014_)
  );
  XOR2X1 _11437_ (
    .A(_05376_),
    .B(_05377_),
    .Y(_04015_)
  );
  NAND2X1 _11438_ (
    .A(_04014_),
    .B(_04015_),
    .Y(_04016_)
  );
  NAND2X1 _11439_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04640_),
    .Y(_04017_)
  );
  NAND2X1 _11440_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04638_),
    .Y(_04018_)
  );
  NAND3X1 _11441_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04642_),
    .C(_05381_),
    .Y(_04019_)
  );
  XNOR2X1 _11442_ (
    .A(_05383_),
    .B(_05385_),
    .Y(_04020_)
  );
  NOR2X1 _11443_ (
    .A(_04019_),
    .B(_04020_),
    .Y(_04021_)
  );
  INVX1 _11444_ (
    .A(_04021_),
    .Y(_04022_)
  );
  XNOR2X1 _11445_ (
    .A(_05364_),
    .B(_05389_),
    .Y(_04023_)
  );
  OR2X1 _11446_ (
    .A(_04022_),
    .B(_04023_),
    .Y(_04024_)
  );
  XNOR2X1 _11447_ (
    .A(_05390_),
    .B(_05391_),
    .Y(_04025_)
  );
  NOR2X1 _11448_ (
    .A(_04024_),
    .B(_04025_),
    .Y(_04026_)
  );
  XOR2X1 _11449_ (
    .A(_05392_),
    .B(_05393_),
    .Y(_04027_)
  );
  NAND2X1 _11450_ (
    .A(_04026_),
    .B(_04027_),
    .Y(_04028_)
  );
  OR2X1 _11451_ (
    .A(_04013_),
    .B(_04028_),
    .Y(_04029_)
  );
  XNOR2X1 _11452_ (
    .A(_04014_),
    .B(_04015_),
    .Y(_04030_)
  );
  OAI21X1 _11453_ (
    .A(_04029_),
    .B(_04030_),
    .C(_04016_),
    .Y(_04031_)
  );
  XOR2X1 _11454_ (
    .A(_05378_),
    .B(_05379_),
    .Y(_04032_)
  );
  AOI21X1 _11455_ (
    .A(_04031_),
    .B(_04032_),
    .C(_05380_),
    .Y(_04033_)
  );
  OAI21X1 _11456_ (
    .A(_05354_),
    .B(_04033_),
    .C(_05353_),
    .Y(_04034_)
  );
  AOI21X1 _11457_ (
    .A(_05320_),
    .B(_04034_),
    .C(_05319_),
    .Y(_04035_)
  );
  OAI21X1 _11458_ (
    .A(_05284_),
    .B(_04035_),
    .C(_05282_),
    .Y(_04036_)
  );
  XOR2X1 _11459_ (
    .A(_05242_),
    .B(_05243_),
    .Y(_04037_)
  );
  AOI21X1 _11460_ (
    .A(_04036_),
    .B(_04037_),
    .C(_05244_),
    .Y(_04038_)
  );
  OAI21X1 _11461_ (
    .A(_05201_),
    .B(_04038_),
    .C(_05199_),
    .Y(_04039_)
  );
  AOI21X1 _11462_ (
    .A(_05158_),
    .B(_04039_),
    .C(_05157_),
    .Y(_04040_)
  );
  OAI21X1 _11463_ (
    .A(_05109_),
    .B(_04040_),
    .C(_05108_),
    .Y(_04041_)
  );
  XOR2X1 _11464_ (
    .A(_05062_),
    .B(_05063_),
    .Y(_04042_)
  );
  AOI21X1 _11465_ (
    .A(_04041_),
    .B(_04042_),
    .C(_05064_),
    .Y(_04043_)
  );
  OAI21X1 _11466_ (
    .A(_05021_),
    .B(_04043_),
    .C(_05019_),
    .Y(_04044_)
  );
  AOI21X1 _11467_ (
    .A(_04976_),
    .B(_04044_),
    .C(_04975_),
    .Y(_04045_)
  );
  OAI21X1 _11468_ (
    .A(_04932_),
    .B(_04045_),
    .C(_04930_),
    .Y(_04046_)
  );
  AOI21X1 _11469_ (
    .A(_04886_),
    .B(_04046_),
    .C(_04885_),
    .Y(_04047_)
  );
  OAI21X1 _11470_ (
    .A(_04842_),
    .B(_04047_),
    .C(_04840_),
    .Y(_04048_)
  );
  XOR2X1 _11471_ (
    .A(_04759_),
    .B(_04794_),
    .Y(_04049_)
  );
  AOI21X1 _11472_ (
    .A(_04048_),
    .B(_04049_),
    .C(_04795_),
    .Y(_04050_)
  );
  OAI21X1 _11473_ (
    .A(_04742_),
    .B(_04754_),
    .C(_04756_),
    .Y(_04051_)
  );
  OAI21X1 _11474_ (
    .A(_04725_),
    .B(_04750_),
    .C(_04752_),
    .Y(_04052_)
  );
  OAI21X1 _11475_ (
    .A(_04734_),
    .B(_04753_),
    .C(_04732_),
    .Y(_04053_)
  );
  NOR2X1 _11476_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04693_),
    .Y(_04054_)
  );
  OAI21X1 _11477_ (
    .A(_04685_),
    .B(_04688_),
    .C(_04643_),
    .Y(_04055_)
  );
  INVX1 _11478_ (
    .A(_04055_),
    .Y(_04056_)
  );
  AOI21X1 _11479_ (
    .A(_04747_),
    .B(_04056_),
    .C(_04054_),
    .Y(_04057_)
  );
  OAI21X1 _11480_ (
    .A(_04749_),
    .B(_04057_),
    .C(_04747_),
    .Y(_04058_)
  );
  XOR2X1 _11481_ (
    .A(_04733_),
    .B(_04058_),
    .Y(_04059_)
  );
  XNOR2X1 _11482_ (
    .A(_04724_),
    .B(_04059_),
    .Y(_04060_)
  );
  XNOR2X1 _11483_ (
    .A(_04053_),
    .B(_04060_),
    .Y(_04061_)
  );
  XNOR2X1 _11484_ (
    .A(_04052_),
    .B(_04061_),
    .Y(_04062_)
  );
  XNOR2X1 _11485_ (
    .A(_04051_),
    .B(_04062_),
    .Y(_04063_)
  );
  XNOR2X1 _11486_ (
    .A(_04758_),
    .B(_04063_),
    .Y(_04064_)
  );
  XNOR2X1 _11487_ (
    .A(_04050_),
    .B(_04064_),
    .Y(_04065_)
  );
  OAI21X1 _11488_ (
    .A( multiplier_0.cycle_0_ ),
    .B( multiplier_0.sign_sel ),
    .C(_04065_),
    .Y(_04066_)
  );
  XNOR2X1 _11489_ (
    .A(_04618_),
    .B(_04066_),
    .Y(_04067_)
  );
  INVX1 _11490_ (
    .A(_04067_),
    .Y(_04068_)
  );
  XNOR2X1 _11491_ (
    .A(_04048_),
    .B(_04049_),
    .Y(_04069_)
  );
  NAND2X1 _11492_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04069_),
    .Y(_04070_)
  );
  NOR2X1 _11493_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04065_),
    .Y(_04071_)
  );
  NOR2X1 _11494_ (
    .A(_04635_),
    .B(_04071_),
    .Y(_04072_)
  );
  INVX1 _11495_ (
    .A(_04072_),
    .Y(_04073_)
  );
  NAND2X1 _11496_ (
    .A(_04070_),
    .B(_04072_),
    .Y(_04074_)
  );
  NAND3X1 _11497_ (
    .A( multiplier_0.reshi_14_ ),
    .B(_04070_),
    .C(_04072_),
    .Y(_04075_)
  );
  XOR2X1 _11498_ (
    .A( multiplier_0.reshi_14_ ),
    .B(_04074_),
    .Y(_04076_)
  );
  XNOR2X1 _11499_ (
    .A(_04841_),
    .B(_04047_),
    .Y(_04077_)
  );
  NOR2X1 _11500_ (
    .A(_04589_),
    .B(_04077_),
    .Y(_04078_)
  );
  NOR2X1 _11501_ (
    .A(_04073_),
    .B(_04078_),
    .Y(_04079_)
  );
  OR2X1 _11502_ (
    .A( multiplier_0.reshi_13_ ),
    .B(_04079_),
    .Y(_04080_)
  );
  NAND2X1 _11503_ (
    .A( multiplier_0.reshi_13_ ),
    .B(_04079_),
    .Y(_04081_)
  );
  INVX1 _11504_ (
    .A(_04081_),
    .Y(_04082_)
  );
  XNOR2X1 _11505_ (
    .A(_04886_),
    .B(_04046_),
    .Y(_04083_)
  );
  AOI21X1 _11506_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04083_),
    .C(_04073_),
    .Y(_04084_)
  );
  NAND2X1 _11507_ (
    .A( multiplier_0.reshi_12_ ),
    .B(_04084_),
    .Y(_04085_)
  );
  XNOR2X1 _11508_ (
    .A( multiplier_0.reshi_12_ ),
    .B(_04084_),
    .Y(_04086_)
  );
  XNOR2X1 _11509_ (
    .A(_04931_),
    .B(_04045_),
    .Y(_04087_)
  );
  NOR2X1 _11510_ (
    .A(_04589_),
    .B(_04087_),
    .Y(_04088_)
  );
  NOR2X1 _11511_ (
    .A(_04073_),
    .B(_04088_),
    .Y(_04089_)
  );
  AND2X1 _11512_ (
    .A( multiplier_0.reshi_11_ ),
    .B(_04089_),
    .Y(_04090_)
  );
  XNOR2X1 _11513_ (
    .A( multiplier_0.reshi_11_ ),
    .B(_04089_),
    .Y(_04091_)
  );
  INVX1 _11514_ (
    .A(_04091_),
    .Y(_04092_)
  );
  XNOR2X1 _11515_ (
    .A(_04976_),
    .B(_04044_),
    .Y(_04093_)
  );
  NAND2X1 _11516_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04093_),
    .Y(_04094_)
  );
  NAND2X1 _11517_ (
    .A(_04072_),
    .B(_04094_),
    .Y(_04095_)
  );
  NAND3X1 _11518_ (
    .A( multiplier_0.reshi_10_ ),
    .B(_04072_),
    .C(_04094_),
    .Y(_04096_)
  );
  XOR2X1 _11519_ (
    .A( multiplier_0.reshi_10_ ),
    .B(_04095_),
    .Y(_04097_)
  );
  XNOR2X1 _11520_ (
    .A(_05021_),
    .B(_04043_),
    .Y(_04098_)
  );
  NAND2X1 _11521_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04098_),
    .Y(_04099_)
  );
  AND2X1 _11522_ (
    .A(_04072_),
    .B(_04099_),
    .Y(_04100_)
  );
  NOR2X1 _11523_ (
    .A( multiplier_0.reshi_9_ ),
    .B(_04100_),
    .Y(_04101_)
  );
  OR2X1 _11524_ (
    .A( multiplier_0.reshi_9_ ),
    .B(_04100_),
    .Y(_04102_)
  );
  AND2X1 _11525_ (
    .A( multiplier_0.reshi_9_ ),
    .B(_04100_),
    .Y(_04103_)
  );
  XNOR2X1 _11526_ (
    .A(_04041_),
    .B(_04042_),
    .Y(_04104_)
  );
  NAND2X1 _11527_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04104_),
    .Y(_04105_)
  );
  NAND2X1 _11528_ (
    .A(_04072_),
    .B(_04105_),
    .Y(_04106_)
  );
  NAND3X1 _11529_ (
    .A( multiplier_0.reshi_8_ ),
    .B(_04072_),
    .C(_04105_),
    .Y(_04107_)
  );
  AOI21X1 _11530_ (
    .A(_04072_),
    .B(_04105_),
    .C( multiplier_0.reshi_8_ ),
    .Y(_04108_)
  );
  XOR2X1 _11531_ (
    .A( multiplier_0.reshi_8_ ),
    .B(_04106_),
    .Y(_04109_)
  );
  XNOR2X1 _11532_ (
    .A(_05110_),
    .B(_04040_),
    .Y(_04110_)
  );
  NOR2X1 _11533_ (
    .A(_04589_),
    .B(_04110_),
    .Y(_04111_)
  );
  NOR2X1 _11534_ (
    .A(_04071_),
    .B(_04111_),
    .Y(_04112_)
  );
  NOR3X1 _11535_ (
    .A(_04617_),
    .B(_04071_),
    .C(_04111_),
    .Y(_04113_)
  );
  NOR2X1 _11536_ (
    .A( multiplier_0.reshi_7_ ),
    .B(_04112_),
    .Y(_04114_)
  );
  OAI21X1 _11537_ (
    .A(_04071_),
    .B(_04111_),
    .C(_04617_),
    .Y(_04115_)
  );
  NOR2X1 _11538_ (
    .A(_04113_),
    .B(_04114_),
    .Y(_04116_)
  );
  XNOR2X1 _11539_ (
    .A(_05158_),
    .B(_04039_),
    .Y(_04117_)
  );
  MUX2X1 _11540_ (
    .A(_04069_),
    .B(_04117_),
    .S(_04589_),
    .Y(_04118_)
  );
  NAND2X1 _11541_ (
    .A( multiplier_0.reshi_6_ ),
    .B(_04118_),
    .Y(_04119_)
  );
  XNOR2X1 _11542_ (
    .A( multiplier_0.reshi_6_ ),
    .B(_04118_),
    .Y(_04120_)
  );
  XNOR2X1 _11543_ (
    .A(_05201_),
    .B(_04038_),
    .Y(_04121_)
  );
  NAND2X1 _11544_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04121_),
    .Y(_04122_)
  );
  OAI21X1 _11545_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04077_),
    .C(_04122_),
    .Y(_04123_)
  );
  NOR2X1 _11546_ (
    .A(_04616_),
    .B(_04123_),
    .Y(_04124_)
  );
  XNOR2X1 _11547_ (
    .A(_04036_),
    .B(_04037_),
    .Y(_04125_)
  );
  MUX2X1 _11548_ (
    .A(_04083_),
    .B(_04125_),
    .S(_04589_),
    .Y(_04126_)
  );
  NAND2X1 _11549_ (
    .A( multiplier_0.reshi_4_ ),
    .B(_04126_),
    .Y(_04127_)
  );
  XNOR2X1 _11550_ (
    .A( multiplier_0.reshi_4_ ),
    .B(_04126_),
    .Y(_04128_)
  );
  XNOR2X1 _11551_ (
    .A(_05283_),
    .B(_04035_),
    .Y(_04129_)
  );
  MUX2X1 _11552_ (
    .A(_04087_),
    .B(_04129_),
    .S(_04589_),
    .Y(_04130_)
  );
  NOR2X1 _11553_ (
    .A(_04615_),
    .B(_04130_),
    .Y(_04131_)
  );
  XNOR2X1 _11554_ (
    .A(_05320_),
    .B(_04034_),
    .Y(_04132_)
  );
  MUX2X1 _11555_ (
    .A(_04093_),
    .B(_04132_),
    .S(_04589_),
    .Y(_04133_)
  );
  NAND2X1 _11556_ (
    .A( multiplier_0.reshi_2_ ),
    .B(_04133_),
    .Y(_04134_)
  );
  XNOR2X1 _11557_ (
    .A( multiplier_0.reshi_2_ ),
    .B(_04133_),
    .Y(_04135_)
  );
  XNOR2X1 _11558_ (
    .A(_05354_),
    .B(_04033_),
    .Y(_04136_)
  );
  MUX2X1 _11559_ (
    .A(_04098_),
    .B(_04136_),
    .S(_04589_),
    .Y(_04137_)
  );
  AND2X1 _11560_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_04137_),
    .Y(_04138_)
  );
  XNOR2X1 _11561_ (
    .A(_04031_),
    .B(_04032_),
    .Y(_04139_)
  );
  MUX2X1 _11562_ (
    .A(_04104_),
    .B(_04139_),
    .S(_04589_),
    .Y(_04140_)
  );
  NAND2X1 _11563_ (
    .A( multiplier_0.reshi_0_ ),
    .B(_04140_),
    .Y(_04141_)
  );
  XNOR2X1 _11564_ (
    .A(_04029_),
    .B(_04030_),
    .Y(_04142_)
  );
  NAND2X1 _11565_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04142_),
    .Y(_04143_)
  );
  OAI21X1 _11566_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04110_),
    .C(_04143_),
    .Y(_04144_)
  );
  NOR2X1 _11567_ (
    .A(_04614_),
    .B(_04144_),
    .Y(_04145_)
  );
  XNOR2X1 _11568_ (
    .A(_04013_),
    .B(_04028_),
    .Y(_04146_)
  );
  AOI21X1 _11569_ (
    .A(_05394_),
    .B(_04146_),
    .C(_04014_),
    .Y(_04147_)
  );
  NAND2X1 _11570_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04147_),
    .Y(_04148_)
  );
  OAI21X1 _11571_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04117_),
    .C(_04148_),
    .Y(_04149_)
  );
  NAND2X1 _11572_ (
    .A( multiplier_0.reslo_14_ ),
    .B(_04149_),
    .Y(_04150_)
  );
  XNOR2X1 _11573_ (
    .A( multiplier_0.reslo_14_ ),
    .B(_04149_),
    .Y(_04151_)
  );
  XNOR2X1 _11574_ (
    .A(_04026_),
    .B(_04027_),
    .Y(_04152_)
  );
  MUX2X1 _11575_ (
    .A(_04121_),
    .B(_04152_),
    .S(_04589_),
    .Y(_04153_)
  );
  AND2X1 _11576_ (
    .A( multiplier_0.reslo_13_ ),
    .B(_04153_),
    .Y(_04154_)
  );
  XOR2X1 _11577_ (
    .A(_04024_),
    .B(_04025_),
    .Y(_04155_)
  );
  NAND2X1 _11578_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04155_),
    .Y(_04156_)
  );
  OAI21X1 _11579_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04125_),
    .C(_04156_),
    .Y(_04157_)
  );
  NAND2X1 _11580_ (
    .A( multiplier_0.reslo_12_ ),
    .B(_04157_),
    .Y(_04158_)
  );
  XNOR2X1 _11581_ (
    .A( multiplier_0.reslo_12_ ),
    .B(_04157_),
    .Y(_04159_)
  );
  XNOR2X1 _11582_ (
    .A(_04021_),
    .B(_04023_),
    .Y(_04160_)
  );
  MUX2X1 _11583_ (
    .A(_04129_),
    .B(_04160_),
    .S(_04589_),
    .Y(_04161_)
  );
  NOR2X1 _11584_ (
    .A(_04612_),
    .B(_04161_),
    .Y(_04162_)
  );
  XNOR2X1 _11585_ (
    .A( multiplier_0.reslo_11_ ),
    .B(_04161_),
    .Y(_04163_)
  );
  XOR2X1 _11586_ (
    .A(_04019_),
    .B(_04020_),
    .Y(_04164_)
  );
  NAND2X1 _11587_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04164_),
    .Y(_04165_)
  );
  OAI21X1 _11588_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04132_),
    .C(_04165_),
    .Y(_04166_)
  );
  NAND2X1 _11589_ (
    .A( multiplier_0.reslo_10_ ),
    .B(_04166_),
    .Y(_04167_)
  );
  XNOR2X1 _11590_ (
    .A( multiplier_0.reslo_10_ ),
    .B(_04166_),
    .Y(_04168_)
  );
  OAI21X1 _11591_ (
    .A(_04596_),
    .B(_04641_),
    .C(_04018_),
    .Y(_04169_)
  );
  AND2X1 _11592_ (
    .A(_04019_),
    .B(_04169_),
    .Y(_04170_)
  );
  NAND2X1 _11593_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04170_),
    .Y(_04171_)
  );
  OAI21X1 _11594_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04136_),
    .C(_04171_),
    .Y(_04172_)
  );
  AND2X1 _11595_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_04172_),
    .Y(_04173_)
  );
  NAND2X1 _11596_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_04172_),
    .Y(_04174_)
  );
  OR2X1 _11597_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_04172_),
    .Y(_04175_)
  );
  NAND2X1 _11598_ (
    .A(_04174_),
    .B(_04175_),
    .Y(_04176_)
  );
  AOI21X1 _11599_ (
    .A( multiplier_0.op2_8_ ),
    .B( multiplier_0.op1_0_ ),
    .C(_04589_),
    .Y(_04177_)
  );
  AOI21X1 _11600_ (
    .A(_04589_),
    .B(_04139_),
    .C(_04177_),
    .Y(_04178_)
  );
  NAND2X1 _11601_ (
    .A( multiplier_0.reslo_8_ ),
    .B(_04178_),
    .Y(_04179_)
  );
  NOR2X1 _11602_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04142_),
    .Y(_04180_)
  );
  AND2X1 _11603_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_04180_),
    .Y(_04181_)
  );
  NAND2X1 _11604_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_04180_),
    .Y(_04182_)
  );
  OR2X1 _11605_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_04180_),
    .Y(_04183_)
  );
  NAND2X1 _11606_ (
    .A(_04182_),
    .B(_04183_),
    .Y(_04184_)
  );
  NAND2X1 _11607_ (
    .A(_04589_),
    .B(_04147_),
    .Y(_04185_)
  );
  NAND3X1 _11608_ (
    .A(_04589_),
    .B( multiplier_0.reslo_6_ ),
    .C(_04147_),
    .Y(_04186_)
  );
  AOI21X1 _11609_ (
    .A(_04589_),
    .B(_04147_),
    .C( multiplier_0.reslo_6_ ),
    .Y(_04187_)
  );
  XNOR2X1 _11610_ (
    .A( multiplier_0.reslo_6_ ),
    .B(_04185_),
    .Y(_04188_)
  );
  NOR2X1 _11611_ (
    .A( multiplier_0.cycle_0_ ),
    .B(_04152_),
    .Y(_04189_)
  );
  AND2X1 _11612_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_04189_),
    .Y(_04190_)
  );
  NAND2X1 _11613_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_04189_),
    .Y(_04191_)
  );
  OR2X1 _11614_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_04189_),
    .Y(_04192_)
  );
  NAND2X1 _11615_ (
    .A(_04191_),
    .B(_04192_),
    .Y(_04193_)
  );
  NAND2X1 _11616_ (
    .A(_04589_),
    .B(_04155_),
    .Y(_04194_)
  );
  NAND3X1 _11617_ (
    .A(_04589_),
    .B( multiplier_0.reslo_4_ ),
    .C(_04155_),
    .Y(_04195_)
  );
  NAND2X1 _11618_ (
    .A(_04589_),
    .B(_04160_),
    .Y(_04196_)
  );
  NAND3X1 _11619_ (
    .A(_04589_),
    .B( multiplier_0.reslo_3_ ),
    .C(_04160_),
    .Y(_04197_)
  );
  AOI21X1 _11620_ (
    .A(_04589_),
    .B(_04160_),
    .C( multiplier_0.reslo_3_ ),
    .Y(_04198_)
  );
  XNOR2X1 _11621_ (
    .A( multiplier_0.reslo_3_ ),
    .B(_04196_),
    .Y(_04199_)
  );
  NAND2X1 _11622_ (
    .A(_04589_),
    .B(_04164_),
    .Y(_04200_)
  );
  NOR2X1 _11623_ (
    .A(_04598_),
    .B(_04200_),
    .Y(_04201_)
  );
  XNOR2X1 _11624_ (
    .A( multiplier_0.reslo_2_ ),
    .B(_04200_),
    .Y(_04202_)
  );
  NAND2X1 _11625_ (
    .A(_04589_),
    .B(_04170_),
    .Y(_04203_)
  );
  NAND3X1 _11626_ (
    .A(_04589_),
    .B( multiplier_0.reslo_1_ ),
    .C(_04170_),
    .Y(_04204_)
  );
  NAND3X1 _11627_ (
    .A( multiplier_0.reslo_0_ ),
    .B( multiplier_0.op1_0_ ),
    .C(_04640_),
    .Y(_04205_)
  );
  AOI21X1 _11628_ (
    .A(_04589_),
    .B(_04170_),
    .C( multiplier_0.reslo_1_ ),
    .Y(_04206_)
  );
  XNOR2X1 _11629_ (
    .A( multiplier_0.reslo_1_ ),
    .B(_04203_),
    .Y(_04207_)
  );
  OAI21X1 _11630_ (
    .A(_04205_),
    .B(_04206_),
    .C(_04204_),
    .Y(_04208_)
  );
  AOI21X1 _11631_ (
    .A(_04202_),
    .B(_04208_),
    .C(_04201_),
    .Y(_04209_)
  );
  OAI21X1 _11632_ (
    .A(_04198_),
    .B(_04209_),
    .C(_04197_),
    .Y(_04210_)
  );
  INVX1 _11633_ (
    .A(_04210_),
    .Y(_04211_)
  );
  XOR2X1 _11634_ (
    .A( multiplier_0.reslo_4_ ),
    .B(_04194_),
    .Y(_04212_)
  );
  OAI21X1 _11635_ (
    .A(_04211_),
    .B(_04212_),
    .C(_04195_),
    .Y(_04213_)
  );
  AOI21X1 _11636_ (
    .A(_04192_),
    .B(_04213_),
    .C(_04190_),
    .Y(_04214_)
  );
  OAI21X1 _11637_ (
    .A(_04187_),
    .B(_04214_),
    .C(_04186_),
    .Y(_04215_)
  );
  AOI21X1 _11638_ (
    .A(_04183_),
    .B(_04215_),
    .C(_04181_),
    .Y(_04216_)
  );
  XNOR2X1 _11639_ (
    .A( multiplier_0.reslo_8_ ),
    .B(_04178_),
    .Y(_04217_)
  );
  OAI21X1 _11640_ (
    .A(_04216_),
    .B(_04217_),
    .C(_04179_),
    .Y(_04218_)
  );
  AOI21X1 _11641_ (
    .A(_04175_),
    .B(_04218_),
    .C(_04173_),
    .Y(_04219_)
  );
  OAI21X1 _11642_ (
    .A(_04168_),
    .B(_04219_),
    .C(_04167_),
    .Y(_04220_)
  );
  AOI21X1 _11643_ (
    .A(_04163_),
    .B(_04220_),
    .C(_04162_),
    .Y(_04221_)
  );
  OAI21X1 _11644_ (
    .A(_04159_),
    .B(_04221_),
    .C(_04158_),
    .Y(_04222_)
  );
  XOR2X1 _11645_ (
    .A( multiplier_0.reslo_13_ ),
    .B(_04153_),
    .Y(_04223_)
  );
  AOI21X1 _11646_ (
    .A(_04222_),
    .B(_04223_),
    .C(_04154_),
    .Y(_04224_)
  );
  OAI21X1 _11647_ (
    .A(_04151_),
    .B(_04224_),
    .C(_04150_),
    .Y(_04225_)
  );
  XNOR2X1 _11648_ (
    .A( multiplier_0.reslo_15_ ),
    .B(_04144_),
    .Y(_04226_)
  );
  AOI21X1 _11649_ (
    .A(_04225_),
    .B(_04226_),
    .C(_04145_),
    .Y(_04227_)
  );
  XNOR2X1 _11650_ (
    .A( multiplier_0.reshi_0_ ),
    .B(_04140_),
    .Y(_04228_)
  );
  OAI21X1 _11651_ (
    .A(_04227_),
    .B(_04228_),
    .C(_04141_),
    .Y(_04229_)
  );
  XOR2X1 _11652_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_04137_),
    .Y(_04230_)
  );
  AOI21X1 _11653_ (
    .A(_04229_),
    .B(_04230_),
    .C(_04138_),
    .Y(_04231_)
  );
  OAI21X1 _11654_ (
    .A(_04135_),
    .B(_04231_),
    .C(_04134_),
    .Y(_04232_)
  );
  XNOR2X1 _11655_ (
    .A( multiplier_0.reshi_3_ ),
    .B(_04130_),
    .Y(_04233_)
  );
  AOI21X1 _11656_ (
    .A(_04232_),
    .B(_04233_),
    .C(_04131_),
    .Y(_04234_)
  );
  OAI21X1 _11657_ (
    .A(_04128_),
    .B(_04234_),
    .C(_04127_),
    .Y(_04235_)
  );
  XNOR2X1 _11658_ (
    .A( multiplier_0.reshi_5_ ),
    .B(_04123_),
    .Y(_04236_)
  );
  AOI21X1 _11659_ (
    .A(_04235_),
    .B(_04236_),
    .C(_04124_),
    .Y(_04237_)
  );
  OAI21X1 _11660_ (
    .A(_04120_),
    .B(_04237_),
    .C(_04119_),
    .Y(_04238_)
  );
  AOI21X1 _11661_ (
    .A(_04115_),
    .B(_04238_),
    .C(_04113_),
    .Y(_04239_)
  );
  OAI21X1 _11662_ (
    .A(_04108_),
    .B(_04239_),
    .C(_04107_),
    .Y(_04240_)
  );
  AOI21X1 _11663_ (
    .A(_04102_),
    .B(_04240_),
    .C(_04103_),
    .Y(_04241_)
  );
  OAI21X1 _11664_ (
    .A(_04097_),
    .B(_04241_),
    .C(_04096_),
    .Y(_04242_)
  );
  AOI21X1 _11665_ (
    .A(_04092_),
    .B(_04242_),
    .C(_04090_),
    .Y(_04243_)
  );
  OAI21X1 _11666_ (
    .A(_04086_),
    .B(_04243_),
    .C(_04085_),
    .Y(_04244_)
  );
  AOI21X1 _11667_ (
    .A(_04080_),
    .B(_04244_),
    .C(_04082_),
    .Y(_04245_)
  );
  OAI21X1 _11668_ (
    .A(_04076_),
    .B(_04245_),
    .C(_04075_),
    .Y(_04246_)
  );
  OAI21X1 _11669_ (
    .A(_04618_),
    .B(_04066_),
    .C(_04619_),
    .Y(_04247_)
  );
  AOI21X1 _11670_ (
    .A(_04068_),
    .B(_04246_),
    .C(_04247_),
    .Y(_04248_)
  );
  NOR2X1 _11671_ (
    .A( multiplier_0.sign_sel ),
    .B(_04248_),
    .Y(_04249_)
  );
  XNOR2X1 _11672_ (
    .A(_04067_),
    .B(_04246_),
    .Y(_04250_)
  );
  AND2X1 _11673_ (
    .A( multiplier_0.sign_sel ),
    .B(_04250_),
    .Y(_04251_)
  );
  AOI21X1 _11674_ (
    .A( multiplier_0.sign_sel ),
    .B(_04250_),
    .C(_04588_),
    .Y(_04252_)
  );
  NOR3X1 _11675_ (
    .A(_04588_),
    .B(_04249_),
    .C(_04251_),
    .Y(_04253_)
  );
  NAND2X1 _11676_ (
    .A(_05635_),
    .B(_05634_),
    .Y(_04254_)
  );
  NAND2X1 _11677_ (
    .A(_04620_),
    .B(_04630_),
    .Y(_04255_)
  );
  NAND3X1 _11678_ (
    .A(_05630_),
    .B(_04620_),
    .C(_04630_),
    .Y(_04256_)
  );
  NOR2X1 _11679_ (
    .A(_04254_),
    .B(_04256_),
    .Y(_04257_)
  );
  OAI21X1 _11680_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.sumext_0_ ),
    .C(_04257_),
    .Y(_04258_)
  );
  XNOR2X1 _11681_ (
    .A(_04227_),
    .B(_04228_),
    .Y(_04259_)
  );
  OR2X1 _11682_ (
    .A(_05630_),
    .B(_04254_),
    .Y(_04260_)
  );
  NOR2X1 _11683_ (
    .A(_04255_),
    .B(_04260_),
    .Y(_04261_)
  );
  OAI21X1 _11684_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_0_ ),
    .C(_04261_),
    .Y(_04262_)
  );
  AOI21X1 _11685_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04259_),
    .C(_04262_),
    .Y(_04263_)
  );
  NOR2X1 _11686_ (
    .A(_04632_),
    .B(_04256_),
    .Y(_04264_)
  );
  INVX1 _11687_ (
    .A(_04264_),
    .Y(_04265_)
  );
  XOR2X1 _11688_ (
    .A( multiplier_0.reslo_0_ ),
    .B(_04017_),
    .Y(_04266_)
  );
  NAND2X1 _11689_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04266_),
    .Y(_04267_)
  );
  OAI21X1 _11690_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_0_ ),
    .C(_04267_),
    .Y(_04268_)
  );
  NOR2X1 _11691_ (
    .A(_05635_),
    .B(_04255_),
    .Y(_04269_)
  );
  NOR2X1 _11692_ (
    .A(_04633_),
    .B(_04255_),
    .Y(_04270_)
  );
  AOI22X1 _11693_ (
    .A( multiplier_0.op1_0_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_0_ ),
    .Y(_04271_)
  );
  OAI21X1 _11694_ (
    .A(_04265_),
    .B(_04268_),
    .C(_04271_),
    .Y(_04272_)
  );
  NOR2X1 _11695_ (
    .A(_04263_),
    .B(_04272_),
    .Y(_04273_)
  );
  OAI21X1 _11696_ (
    .A(_04253_),
    .B(_04258_),
    .C(_04273_),
    .Y( multiplier_0.per_dout_0_ )
  );
  OAI21X1 _11697_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.sumext_10_ ),
    .C(_04257_),
    .Y(_04274_)
  );
  OR2X1 _11698_ (
    .A(_04252_),
    .B(_04274_),
    .Y(_04275_)
  );
  XNOR2X1 _11699_ (
    .A(_04229_),
    .B(_04230_),
    .Y(_04276_)
  );
  OAI21X1 _11700_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_1_ ),
    .C(_04261_),
    .Y(_04277_)
  );
  AOI21X1 _11701_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04276_),
    .C(_04277_),
    .Y(_04278_)
  );
  XOR2X1 _11702_ (
    .A(_04205_),
    .B(_04207_),
    .Y(_04279_)
  );
  AND2X1 _11703_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04279_),
    .Y(_04280_)
  );
  OAI21X1 _11704_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_1_ ),
    .C(_04264_),
    .Y(_04281_)
  );
  AOI22X1 _11705_ (
    .A( multiplier_0.op1_1_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_1_ ),
    .Y(_04282_)
  );
  OAI21X1 _11706_ (
    .A(_04280_),
    .B(_04281_),
    .C(_04282_),
    .Y(_04283_)
  );
  NOR2X1 _11707_ (
    .A(_04278_),
    .B(_04283_),
    .Y(_04284_)
  );
  OAI21X1 _11708_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04284_),
    .Y( multiplier_0.per_dout_1_ )
  );
  XNOR2X1 _11709_ (
    .A(_04135_),
    .B(_04231_),
    .Y(_04285_)
  );
  OAI21X1 _11710_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_2_ ),
    .C(_04261_),
    .Y(_04286_)
  );
  AOI21X1 _11711_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04285_),
    .C(_04286_),
    .Y(_04287_)
  );
  XNOR2X1 _11712_ (
    .A(_04202_),
    .B(_04208_),
    .Y(_04288_)
  );
  AND2X1 _11713_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04288_),
    .Y(_04289_)
  );
  OAI21X1 _11714_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_2_ ),
    .C(_04264_),
    .Y(_04290_)
  );
  AOI22X1 _11715_ (
    .A( multiplier_0.op1_2_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_2_ ),
    .Y(_04291_)
  );
  OAI21X1 _11716_ (
    .A(_04289_),
    .B(_04290_),
    .C(_04291_),
    .Y(_04292_)
  );
  NOR2X1 _11717_ (
    .A(_04287_),
    .B(_04292_),
    .Y(_04293_)
  );
  OAI21X1 _11718_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04293_),
    .Y( multiplier_0.per_dout_2_ )
  );
  XNOR2X1 _11719_ (
    .A(_04232_),
    .B(_04233_),
    .Y(_04294_)
  );
  OAI21X1 _11720_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_3_ ),
    .C(_04261_),
    .Y(_04295_)
  );
  AOI21X1 _11721_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04294_),
    .C(_04295_),
    .Y(_04296_)
  );
  XNOR2X1 _11722_ (
    .A(_04199_),
    .B(_04209_),
    .Y(_04297_)
  );
  INVX1 _11723_ (
    .A(_04297_),
    .Y(_04298_)
  );
  NOR2X1 _11724_ (
    .A(_04588_),
    .B(_04297_),
    .Y(_04299_)
  );
  OAI21X1 _11725_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_3_ ),
    .C(_04264_),
    .Y(_04300_)
  );
  AOI22X1 _11726_ (
    .A( multiplier_0.op1_3_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_3_ ),
    .Y(_04301_)
  );
  OAI21X1 _11727_ (
    .A(_04299_),
    .B(_04300_),
    .C(_04301_),
    .Y(_04302_)
  );
  NOR2X1 _11728_ (
    .A(_04296_),
    .B(_04302_),
    .Y(_04303_)
  );
  OAI21X1 _11729_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04303_),
    .Y( multiplier_0.per_dout_3_ )
  );
  XNOR2X1 _11730_ (
    .A(_04128_),
    .B(_04234_),
    .Y(_04304_)
  );
  OAI21X1 _11731_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_4_ ),
    .C(_04261_),
    .Y(_04305_)
  );
  AOI21X1 _11732_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04304_),
    .C(_04305_),
    .Y(_04306_)
  );
  XNOR2X1 _11733_ (
    .A(_04210_),
    .B(_04212_),
    .Y(_04307_)
  );
  INVX1 _11734_ (
    .A(_04307_),
    .Y(_04308_)
  );
  NOR2X1 _11735_ (
    .A(_04588_),
    .B(_04307_),
    .Y(_04309_)
  );
  OAI21X1 _11736_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_4_ ),
    .C(_04264_),
    .Y(_04310_)
  );
  AOI22X1 _11737_ (
    .A( multiplier_0.op1_4_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_4_ ),
    .Y(_04311_)
  );
  OAI21X1 _11738_ (
    .A(_04309_),
    .B(_04310_),
    .C(_04311_),
    .Y(_04312_)
  );
  NOR2X1 _11739_ (
    .A(_04306_),
    .B(_04312_),
    .Y(_04313_)
  );
  OAI21X1 _11740_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04313_),
    .Y( multiplier_0.per_dout_4_ )
  );
  XNOR2X1 _11741_ (
    .A(_04235_),
    .B(_04236_),
    .Y(_04314_)
  );
  OAI21X1 _11742_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_5_ ),
    .C(_04261_),
    .Y(_04315_)
  );
  AOI21X1 _11743_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04314_),
    .C(_04315_),
    .Y(_04316_)
  );
  XNOR2X1 _11744_ (
    .A(_04193_),
    .B(_04213_),
    .Y(_04317_)
  );
  INVX1 _11745_ (
    .A(_04317_),
    .Y(_04318_)
  );
  NOR2X1 _11746_ (
    .A(_04588_),
    .B(_04317_),
    .Y(_04319_)
  );
  OAI21X1 _11747_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_5_ ),
    .C(_04264_),
    .Y(_04320_)
  );
  AOI22X1 _11748_ (
    .A( multiplier_0.op1_5_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_5_ ),
    .Y(_04321_)
  );
  OAI21X1 _11749_ (
    .A(_04319_),
    .B(_04320_),
    .C(_04321_),
    .Y(_04322_)
  );
  NOR2X1 _11750_ (
    .A(_04316_),
    .B(_04322_),
    .Y(_04323_)
  );
  OAI21X1 _11751_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04323_),
    .Y( multiplier_0.per_dout_5_ )
  );
  XNOR2X1 _11752_ (
    .A(_04120_),
    .B(_04237_),
    .Y(_04324_)
  );
  OAI21X1 _11753_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_6_ ),
    .C(_04261_),
    .Y(_04325_)
  );
  AOI21X1 _11754_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04324_),
    .C(_04325_),
    .Y(_04326_)
  );
  XOR2X1 _11755_ (
    .A(_04188_),
    .B(_04214_),
    .Y(_04327_)
  );
  AND2X1 _11756_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04327_),
    .Y(_04328_)
  );
  OAI21X1 _11757_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_6_ ),
    .C(_04264_),
    .Y(_04329_)
  );
  AOI22X1 _11758_ (
    .A( multiplier_0.op1_6_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_6_ ),
    .Y(_04330_)
  );
  OAI21X1 _11759_ (
    .A(_04328_),
    .B(_04329_),
    .C(_04330_),
    .Y(_04331_)
  );
  NOR2X1 _11760_ (
    .A(_04326_),
    .B(_04331_),
    .Y(_04332_)
  );
  OAI21X1 _11761_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04332_),
    .Y( multiplier_0.per_dout_6_ )
  );
  XNOR2X1 _11762_ (
    .A(_04116_),
    .B(_04238_),
    .Y(_04333_)
  );
  OAI21X1 _11763_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_7_ ),
    .C(_04261_),
    .Y(_04334_)
  );
  AOI21X1 _11764_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04333_),
    .C(_04334_),
    .Y(_04335_)
  );
  XNOR2X1 _11765_ (
    .A(_04184_),
    .B(_04215_),
    .Y(_04336_)
  );
  INVX1 _11766_ (
    .A(_04336_),
    .Y(_04337_)
  );
  NOR2X1 _11767_ (
    .A(_04588_),
    .B(_04336_),
    .Y(_04338_)
  );
  OAI21X1 _11768_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_7_ ),
    .C(_04264_),
    .Y(_04339_)
  );
  AOI22X1 _11769_ (
    .A( multiplier_0.op1_7_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_7_ ),
    .Y(_04340_)
  );
  OAI21X1 _11770_ (
    .A(_04338_),
    .B(_04339_),
    .C(_04340_),
    .Y(_04341_)
  );
  NOR2X1 _11771_ (
    .A(_04335_),
    .B(_04341_),
    .Y(_04342_)
  );
  OAI21X1 _11772_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04342_),
    .Y( multiplier_0.per_dout_7_ )
  );
  XNOR2X1 _11773_ (
    .A(_04109_),
    .B(_04239_),
    .Y(_04343_)
  );
  OAI21X1 _11774_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_8_ ),
    .C(_04261_),
    .Y(_04344_)
  );
  AOI21X1 _11775_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04343_),
    .C(_04344_),
    .Y(_04345_)
  );
  XNOR2X1 _11776_ (
    .A(_04216_),
    .B(_04217_),
    .Y(_04346_)
  );
  AND2X1 _11777_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04346_),
    .Y(_04347_)
  );
  OAI21X1 _11778_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_8_ ),
    .C(_04264_),
    .Y(_04348_)
  );
  AOI22X1 _11779_ (
    .A( multiplier_0.op1_8_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_8_ ),
    .Y(_04349_)
  );
  OAI21X1 _11780_ (
    .A(_04347_),
    .B(_04348_),
    .C(_04349_),
    .Y(_04350_)
  );
  NOR2X1 _11781_ (
    .A(_04345_),
    .B(_04350_),
    .Y(_04351_)
  );
  OAI21X1 _11782_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04351_),
    .Y( multiplier_0.per_dout_8_ )
  );
  NOR2X1 _11783_ (
    .A(_04101_),
    .B(_04103_),
    .Y(_04352_)
  );
  XNOR2X1 _11784_ (
    .A(_04240_),
    .B(_04352_),
    .Y(_04353_)
  );
  OAI21X1 _11785_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_9_ ),
    .C(_04261_),
    .Y(_04354_)
  );
  AOI21X1 _11786_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04353_),
    .C(_04354_),
    .Y(_04355_)
  );
  XOR2X1 _11787_ (
    .A(_04176_),
    .B(_04218_),
    .Y(_04356_)
  );
  AND2X1 _11788_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04356_),
    .Y(_04357_)
  );
  OAI21X1 _11789_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_9_ ),
    .C(_04264_),
    .Y(_04358_)
  );
  AOI22X1 _11790_ (
    .A( multiplier_0.op1_9_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_9_ ),
    .Y(_04359_)
  );
  OAI21X1 _11791_ (
    .A(_04357_),
    .B(_04358_),
    .C(_04359_),
    .Y(_04360_)
  );
  NOR2X1 _11792_ (
    .A(_04355_),
    .B(_04360_),
    .Y(_04361_)
  );
  OAI21X1 _11793_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04361_),
    .Y( multiplier_0.per_dout_9_ )
  );
  XNOR2X1 _11794_ (
    .A(_04097_),
    .B(_04241_),
    .Y(_04362_)
  );
  OAI21X1 _11795_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_10_ ),
    .C(_04261_),
    .Y(_04363_)
  );
  AOI21X1 _11796_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04362_),
    .C(_04363_),
    .Y(_04364_)
  );
  XNOR2X1 _11797_ (
    .A(_04168_),
    .B(_04219_),
    .Y(_04365_)
  );
  AND2X1 _11798_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04365_),
    .Y(_04366_)
  );
  OAI21X1 _11799_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_10_ ),
    .C(_04264_),
    .Y(_04367_)
  );
  AOI22X1 _11800_ (
    .A( multiplier_0.op1_10_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_10_ ),
    .Y(_04368_)
  );
  OAI21X1 _11801_ (
    .A(_04366_),
    .B(_04367_),
    .C(_04368_),
    .Y(_04369_)
  );
  NOR2X1 _11802_ (
    .A(_04364_),
    .B(_04369_),
    .Y(_04370_)
  );
  OAI21X1 _11803_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04370_),
    .Y( multiplier_0.per_dout_10_ )
  );
  XNOR2X1 _11804_ (
    .A(_04092_),
    .B(_04242_),
    .Y(_04371_)
  );
  OAI21X1 _11805_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_11_ ),
    .C(_04261_),
    .Y(_04372_)
  );
  AOI21X1 _11806_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04371_),
    .C(_04372_),
    .Y(_04373_)
  );
  XNOR2X1 _11807_ (
    .A(_04163_),
    .B(_04220_),
    .Y(_04374_)
  );
  AND2X1 _11808_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04374_),
    .Y(_04375_)
  );
  OAI21X1 _11809_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_11_ ),
    .C(_04264_),
    .Y(_04376_)
  );
  AOI22X1 _11810_ (
    .A( multiplier_0.op1_11_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_11_ ),
    .Y(_04377_)
  );
  OAI21X1 _11811_ (
    .A(_04375_),
    .B(_04376_),
    .C(_04377_),
    .Y(_04378_)
  );
  NOR2X1 _11812_ (
    .A(_04373_),
    .B(_04378_),
    .Y(_04379_)
  );
  OAI21X1 _11813_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04379_),
    .Y( multiplier_0.per_dout_11_ )
  );
  XNOR2X1 _11814_ (
    .A(_04086_),
    .B(_04243_),
    .Y(_04380_)
  );
  OAI21X1 _11815_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_12_ ),
    .C(_04261_),
    .Y(_04381_)
  );
  AOI21X1 _11816_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04380_),
    .C(_04381_),
    .Y(_04382_)
  );
  XNOR2X1 _11817_ (
    .A(_04159_),
    .B(_04221_),
    .Y(_04383_)
  );
  AND2X1 _11818_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04383_),
    .Y(_04384_)
  );
  OAI21X1 _11819_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_12_ ),
    .C(_04264_),
    .Y(_04385_)
  );
  AOI22X1 _11820_ (
    .A( multiplier_0.op1_12_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_12_ ),
    .Y(_04386_)
  );
  OAI21X1 _11821_ (
    .A(_04384_),
    .B(_04385_),
    .C(_04386_),
    .Y(_04387_)
  );
  NOR2X1 _11822_ (
    .A(_04382_),
    .B(_04387_),
    .Y(_04388_)
  );
  OAI21X1 _11823_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04388_),
    .Y( multiplier_0.per_dout_12_ )
  );
  NAND2X1 _11824_ (
    .A(_04080_),
    .B(_04081_),
    .Y(_04389_)
  );
  XOR2X1 _11825_ (
    .A(_04244_),
    .B(_04389_),
    .Y(_04390_)
  );
  OAI21X1 _11826_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_13_ ),
    .C(_04261_),
    .Y(_04391_)
  );
  AOI21X1 _11827_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04390_),
    .C(_04391_),
    .Y(_04392_)
  );
  XNOR2X1 _11828_ (
    .A(_04222_),
    .B(_04223_),
    .Y(_04393_)
  );
  AND2X1 _11829_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04393_),
    .Y(_04394_)
  );
  OAI21X1 _11830_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_13_ ),
    .C(_04264_),
    .Y(_04395_)
  );
  AOI22X1 _11831_ (
    .A( multiplier_0.op1_13_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_13_ ),
    .Y(_04396_)
  );
  OAI21X1 _11832_ (
    .A(_04394_),
    .B(_04395_),
    .C(_04396_),
    .Y(_04397_)
  );
  NOR2X1 _11833_ (
    .A(_04392_),
    .B(_04397_),
    .Y(_04398_)
  );
  OAI21X1 _11834_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04398_),
    .Y( multiplier_0.per_dout_13_ )
  );
  XNOR2X1 _11835_ (
    .A(_04076_),
    .B(_04245_),
    .Y(_04399_)
  );
  OAI21X1 _11836_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_14_ ),
    .C(_04261_),
    .Y(_04400_)
  );
  AOI21X1 _11837_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04399_),
    .C(_04400_),
    .Y(_04401_)
  );
  XNOR2X1 _11838_ (
    .A(_04151_),
    .B(_04224_),
    .Y(_04402_)
  );
  AND2X1 _11839_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04402_),
    .Y(_04403_)
  );
  OAI21X1 _11840_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_14_ ),
    .C(_04264_),
    .Y(_04404_)
  );
  AOI22X1 _11841_ (
    .A( multiplier_0.op1_14_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_14_ ),
    .Y(_04405_)
  );
  OAI21X1 _11842_ (
    .A(_04403_),
    .B(_04404_),
    .C(_04405_),
    .Y(_04406_)
  );
  NOR2X1 _11843_ (
    .A(_04401_),
    .B(_04406_),
    .Y(_04407_)
  );
  OAI21X1 _11844_ (
    .A(_04252_),
    .B(_04274_),
    .C(_04407_),
    .Y( multiplier_0.per_dout_14_ )
  );
  OAI21X1 _11845_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reshi_15_ ),
    .C(_04261_),
    .Y(_04408_)
  );
  INVX1 _11846_ (
    .A(_04408_),
    .Y(_04409_)
  );
  OAI21X1 _11847_ (
    .A(_04588_),
    .B(_04250_),
    .C(_04409_),
    .Y(_04410_)
  );
  XNOR2X1 _11848_ (
    .A(_04225_),
    .B(_04226_),
    .Y(_04411_)
  );
  AND2X1 _11849_ (
    .A( multiplier_0.cycle_1_ ),
    .B(_04411_),
    .Y(_04412_)
  );
  OAI21X1 _11850_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.reslo_15_ ),
    .C(_04264_),
    .Y(_04413_)
  );
  AOI22X1 _11851_ (
    .A( multiplier_0.op1_15_ ),
    .B(_04269_),
    .C(_04270_),
    .D( multiplier_0.op2_15_ ),
    .Y(_04414_)
  );
  OAI21X1 _11852_ (
    .A(_04412_),
    .B(_04413_),
    .C(_04414_),
    .Y(_04415_)
  );
  INVX1 _11853_ (
    .A(_04415_),
    .Y(_04416_)
  );
  NAND3X1 _11854_ (
    .A(_04275_),
    .B(_04410_),
    .C(_04416_),
    .Y( multiplier_0.per_dout_15_ )
  );
  NOR2X1 _11855_ (
    .A(_04593_),
    .B(_05642_),
    .Y(_04417_)
  );
  NAND3X1 _11856_ (
    .A(_05636_),
    .B(_04592_),
    .C(_04417_),
    .Y(_04418_)
  );
  NOR2X1 _11857_ (
    .A(_05641_),
    .B(_05631_),
    .Y(_04419_)
  );
  NOR2X1 _11858_ (
    .A(_04591_),
    .B(_05638_),
    .Y(_04420_)
  );
  NAND3X1 _11859_ (
    .A(_04623_),
    .B(_04419_),
    .C(_04420_),
    .Y(_04421_)
  );
  NOR2X1 _11860_ (
    .A(_04418_),
    .B(_04421_),
    .Y(_04422_)
  );
  OAI21X1 _11861_ (
    .A(_05661_),
    .B(_05660_),
    .C(_04422_),
    .Y(_04423_)
  );
  OR2X1 _11862_ (
    .A(_05635_),
    .B(_04423_),
    .Y(_04424_)
  );
  MUX2X1 _11863_ (
    .A( multiplier_0.acc_sel ),
    .B(_05634_),
    .S(_04424_),
    .Y(_04425_)
  );
  INVX1 _11864_ (
    .A(_04425_),
    .Y(_03945_)
  );
  MUX2X1 _11865_ (
    .A( multiplier_0.sign_sel ),
    .B(_05630_),
    .S(_04424_),
    .Y(_04426_)
  );
  INVX1 _11866_ (
    .A(_04426_),
    .Y(_03946_)
  );
  NOR2X1 _11867_ (
    .A( multiplier_0.cycle_1_ ),
    .B( multiplier_0.cycle_0_ ),
    .Y(_04427_)
  );
  NAND2X1 _11868_ (
    .A(_04588_),
    .B(_04589_),
    .Y(_04428_)
  );
  OR2X1 _11869_ (
    .A(_04633_),
    .B(_04423_),
    .Y(_04429_)
  );
  NAND3X1 _11870_ (
    .A(_04251_),
    .B(_04428_),
    .C(_04429_),
    .Y(_04430_)
  );
  NAND3X1 _11871_ (
    .A( multiplier_0.sumext_0_ ),
    .B(_04427_),
    .C(_04429_),
    .Y(_04431_)
  );
  NAND3X1 _11872_ (
    .A(_04249_),
    .B(_04428_),
    .C(_04429_),
    .Y(_04432_)
  );
  NAND3X1 _11873_ (
    .A(_04430_),
    .B(_04431_),
    .C(_04432_),
    .Y(_03947_)
  );
  NAND3X1 _11874_ (
    .A( multiplier_0.sumext_10_ ),
    .B(_04427_),
    .C(_04429_),
    .Y(_04433_)
  );
  NAND2X1 _11875_ (
    .A(_04430_),
    .B(_04433_),
    .Y(_03948_)
  );
  NOR2X1 _11876_ (
    .A(_04631_),
    .B(_04260_),
    .Y(_04434_)
  );
  INVX1 _11877_ (
    .A(_04434_),
    .Y(_04435_)
  );
  OAI21X1 _11878_ (
    .A( multiplier_0.acc_sel ),
    .B(_04634_),
    .C(_04435_),
    .Y(_04436_)
  );
  INVX1 _11879_ (
    .A(_04436_),
    .Y(_04437_)
  );
  NOR2X1 _11880_ (
    .A(_04428_),
    .B(_04436_),
    .Y(_04438_)
  );
  NAND2X1 _11881_ (
    .A(_04427_),
    .B(_04437_),
    .Y(_04439_)
  );
  AOI21X1 _11882_ (
    .A(_05643_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04440_)
  );
  OAI21X1 _11883_ (
    .A(_04259_),
    .B(_04436_),
    .C(_04440_),
    .Y(_04441_)
  );
  OAI21X1 _11884_ (
    .A( multiplier_0.reshi_0_ ),
    .B(_04439_),
    .C(_04441_),
    .Y(_04442_)
  );
  INVX1 _11885_ (
    .A(_04442_),
    .Y(_03949_)
  );
  AOI21X1 _11886_ (
    .A(_05650_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04443_)
  );
  OAI21X1 _11887_ (
    .A(_04276_),
    .B(_04436_),
    .C(_04443_),
    .Y(_04444_)
  );
  OAI21X1 _11888_ (
    .A( multiplier_0.reshi_1_ ),
    .B(_04439_),
    .C(_04444_),
    .Y(_04445_)
  );
  INVX1 _11889_ (
    .A(_04445_),
    .Y(_03950_)
  );
  AOI21X1 _11890_ (
    .A(_05651_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04446_)
  );
  OAI21X1 _11891_ (
    .A(_04285_),
    .B(_04436_),
    .C(_04446_),
    .Y(_04447_)
  );
  OAI21X1 _11892_ (
    .A( multiplier_0.reshi_2_ ),
    .B(_04439_),
    .C(_04447_),
    .Y(_04448_)
  );
  INVX1 _11893_ (
    .A(_04448_),
    .Y(_03951_)
  );
  AOI21X1 _11894_ (
    .A(_05652_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04449_)
  );
  OAI21X1 _11895_ (
    .A(_04294_),
    .B(_04436_),
    .C(_04449_),
    .Y(_04450_)
  );
  OAI21X1 _11896_ (
    .A( multiplier_0.reshi_3_ ),
    .B(_04439_),
    .C(_04450_),
    .Y(_04451_)
  );
  INVX1 _11897_ (
    .A(_04451_),
    .Y(_03952_)
  );
  AOI21X1 _11898_ (
    .A(_05653_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04452_)
  );
  OAI21X1 _11899_ (
    .A(_04304_),
    .B(_04436_),
    .C(_04452_),
    .Y(_04453_)
  );
  OAI21X1 _11900_ (
    .A( multiplier_0.reshi_4_ ),
    .B(_04439_),
    .C(_04453_),
    .Y(_04454_)
  );
  INVX1 _11901_ (
    .A(_04454_),
    .Y(_03953_)
  );
  AOI21X1 _11902_ (
    .A(_05654_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04455_)
  );
  OAI21X1 _11903_ (
    .A(_04314_),
    .B(_04436_),
    .C(_04455_),
    .Y(_04456_)
  );
  OAI21X1 _11904_ (
    .A( multiplier_0.reshi_5_ ),
    .B(_04439_),
    .C(_04456_),
    .Y(_04457_)
  );
  INVX1 _11905_ (
    .A(_04457_),
    .Y(_03954_)
  );
  AOI21X1 _11906_ (
    .A(_05655_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04458_)
  );
  OAI21X1 _11907_ (
    .A(_04324_),
    .B(_04436_),
    .C(_04458_),
    .Y(_04459_)
  );
  OAI21X1 _11908_ (
    .A( multiplier_0.reshi_6_ ),
    .B(_04439_),
    .C(_04459_),
    .Y(_04460_)
  );
  INVX1 _11909_ (
    .A(_04460_),
    .Y(_03955_)
  );
  AOI21X1 _11910_ (
    .A(_05656_),
    .B(_04434_),
    .C(_04438_),
    .Y(_04461_)
  );
  OAI21X1 _11911_ (
    .A(_04333_),
    .B(_04436_),
    .C(_04461_),
    .Y(_04462_)
  );
  OAI21X1 _11912_ (
    .A( multiplier_0.reshi_7_ ),
    .B(_04439_),
    .C(_04462_),
    .Y(_04463_)
  );
  INVX1 _11913_ (
    .A(_04463_),
    .Y(_03956_)
  );
  AND2X1 _11914_ (
    .A(_05661_),
    .B(_05657_),
    .Y(_04464_)
  );
  NAND2X1 _11915_ (
    .A(_05661_),
    .B(_05657_),
    .Y(_04465_)
  );
  AOI21X1 _11916_ (
    .A(_04434_),
    .B(_04464_),
    .C(_04438_),
    .Y(_04466_)
  );
  OAI21X1 _11917_ (
    .A(_04343_),
    .B(_04436_),
    .C(_04466_),
    .Y(_04467_)
  );
  OAI21X1 _11918_ (
    .A( multiplier_0.reshi_8_ ),
    .B(_04439_),
    .C(_04467_),
    .Y(_04468_)
  );
  INVX1 _11919_ (
    .A(_04468_),
    .Y(_03957_)
  );
  AND2X1 _11920_ (
    .A(_05661_),
    .B(_05658_),
    .Y(_04469_)
  );
  NAND2X1 _11921_ (
    .A(_05661_),
    .B(_05658_),
    .Y(_04470_)
  );
  AOI21X1 _11922_ (
    .A(_04434_),
    .B(_04469_),
    .C(_04438_),
    .Y(_04471_)
  );
  OAI21X1 _11923_ (
    .A(_04353_),
    .B(_04436_),
    .C(_04471_),
    .Y(_04472_)
  );
  OAI21X1 _11924_ (
    .A( multiplier_0.reshi_9_ ),
    .B(_04439_),
    .C(_04472_),
    .Y(_04473_)
  );
  INVX1 _11925_ (
    .A(_04473_),
    .Y(_03958_)
  );
  AND2X1 _11926_ (
    .A(_05661_),
    .B(_05644_),
    .Y(_04474_)
  );
  NAND2X1 _11927_ (
    .A(_05661_),
    .B(_05644_),
    .Y(_04475_)
  );
  AOI21X1 _11928_ (
    .A(_04434_),
    .B(_04474_),
    .C(_04438_),
    .Y(_04476_)
  );
  OAI21X1 _11929_ (
    .A(_04362_),
    .B(_04436_),
    .C(_04476_),
    .Y(_04477_)
  );
  OAI21X1 _11930_ (
    .A( multiplier_0.reshi_10_ ),
    .B(_04439_),
    .C(_04477_),
    .Y(_04478_)
  );
  INVX1 _11931_ (
    .A(_04478_),
    .Y(_03959_)
  );
  AND2X1 _11932_ (
    .A(_05661_),
    .B(_05645_),
    .Y(_04479_)
  );
  NAND2X1 _11933_ (
    .A(_05661_),
    .B(_05645_),
    .Y(_04480_)
  );
  AOI21X1 _11934_ (
    .A(_04434_),
    .B(_04479_),
    .C(_04438_),
    .Y(_04481_)
  );
  OAI21X1 _11935_ (
    .A(_04371_),
    .B(_04436_),
    .C(_04481_),
    .Y(_04482_)
  );
  OAI21X1 _11936_ (
    .A( multiplier_0.reshi_11_ ),
    .B(_04439_),
    .C(_04482_),
    .Y(_04483_)
  );
  INVX1 _11937_ (
    .A(_04483_),
    .Y(_03960_)
  );
  AND2X1 _11938_ (
    .A(_05661_),
    .B(_05646_),
    .Y(_04484_)
  );
  NAND2X1 _11939_ (
    .A(_05661_),
    .B(_05646_),
    .Y(_04485_)
  );
  AOI21X1 _11940_ (
    .A(_04434_),
    .B(_04484_),
    .C(_04438_),
    .Y(_04486_)
  );
  OAI21X1 _11941_ (
    .A(_04380_),
    .B(_04436_),
    .C(_04486_),
    .Y(_04487_)
  );
  OAI21X1 _11942_ (
    .A( multiplier_0.reshi_12_ ),
    .B(_04439_),
    .C(_04487_),
    .Y(_04488_)
  );
  INVX1 _11943_ (
    .A(_04488_),
    .Y(_03961_)
  );
  AND2X1 _11944_ (
    .A(_05661_),
    .B(_05647_),
    .Y(_04489_)
  );
  NAND2X1 _11945_ (
    .A(_05661_),
    .B(_05647_),
    .Y(_04490_)
  );
  AOI21X1 _11946_ (
    .A(_04434_),
    .B(_04489_),
    .C(_04438_),
    .Y(_04491_)
  );
  OAI21X1 _11947_ (
    .A(_04390_),
    .B(_04436_),
    .C(_04491_),
    .Y(_04492_)
  );
  OAI21X1 _11948_ (
    .A( multiplier_0.reshi_13_ ),
    .B(_04439_),
    .C(_04492_),
    .Y(_04493_)
  );
  INVX1 _11949_ (
    .A(_04493_),
    .Y(_03962_)
  );
  AND2X1 _11950_ (
    .A(_05661_),
    .B(_05648_),
    .Y(_04494_)
  );
  NAND2X1 _11951_ (
    .A(_05661_),
    .B(_05648_),
    .Y(_04495_)
  );
  AOI21X1 _11952_ (
    .A(_04434_),
    .B(_04494_),
    .C(_04438_),
    .Y(_04496_)
  );
  OAI21X1 _11953_ (
    .A(_04399_),
    .B(_04436_),
    .C(_04496_),
    .Y(_04497_)
  );
  OAI21X1 _11954_ (
    .A( multiplier_0.reshi_14_ ),
    .B(_04439_),
    .C(_04497_),
    .Y(_04498_)
  );
  INVX1 _11955_ (
    .A(_04498_),
    .Y(_03963_)
  );
  NAND2X1 _11956_ (
    .A(_05661_),
    .B(_05649_),
    .Y(_04499_)
  );
  OAI21X1 _11957_ (
    .A(_04435_),
    .B(_04499_),
    .C(_04439_),
    .Y(_04500_)
  );
  AOI21X1 _11958_ (
    .A(_04250_),
    .B(_04437_),
    .C(_04500_),
    .Y(_04501_)
  );
  AOI21X1 _11959_ (
    .A(_04618_),
    .B(_04438_),
    .C(_04501_),
    .Y(_03964_)
  );
  NAND3X1 _11960_ (
    .A(_05635_),
    .B(_04590_),
    .C(_05630_),
    .Y(_04502_)
  );
  NOR2X1 _11961_ (
    .A(_04631_),
    .B(_04502_),
    .Y(_04503_)
  );
  INVX1 _11962_ (
    .A(_04503_),
    .Y(_04504_)
  );
  OAI21X1 _11963_ (
    .A( multiplier_0.acc_sel ),
    .B(_04634_),
    .C(_04504_),
    .Y(_04505_)
  );
  NOR2X1 _11964_ (
    .A(_04428_),
    .B(_04505_),
    .Y(_04506_)
  );
  OR2X1 _11965_ (
    .A(_04428_),
    .B(_04505_),
    .Y(_04507_)
  );
  NOR2X1 _11966_ (
    .A(_04266_),
    .B(_04505_),
    .Y(_04508_)
  );
  AOI21X1 _11967_ (
    .A(_05643_),
    .B(_04503_),
    .C(_04508_),
    .Y(_04509_)
  );
  NAND2X1 _11968_ (
    .A( multiplier_0.reslo_0_ ),
    .B(_04506_),
    .Y(_04510_)
  );
  OAI21X1 _11969_ (
    .A(_04506_),
    .B(_04509_),
    .C(_04510_),
    .Y(_03965_)
  );
  NOR2X1 _11970_ (
    .A(_04279_),
    .B(_04505_),
    .Y(_04511_)
  );
  AOI21X1 _11971_ (
    .A(_05650_),
    .B(_04503_),
    .C(_04511_),
    .Y(_04512_)
  );
  NAND2X1 _11972_ (
    .A( multiplier_0.reslo_1_ ),
    .B(_04506_),
    .Y(_04513_)
  );
  OAI21X1 _11973_ (
    .A(_04506_),
    .B(_04512_),
    .C(_04513_),
    .Y(_03966_)
  );
  NAND2X1 _11974_ (
    .A(_05651_),
    .B(_04503_),
    .Y(_04514_)
  );
  OAI21X1 _11975_ (
    .A(_04288_),
    .B(_04505_),
    .C(_04514_),
    .Y(_04515_)
  );
  OAI21X1 _11976_ (
    .A(_04428_),
    .B(_04505_),
    .C(_04515_),
    .Y(_04516_)
  );
  OAI21X1 _11977_ (
    .A(_04598_),
    .B(_04507_),
    .C(_04516_),
    .Y(_03967_)
  );
  AOI21X1 _11978_ (
    .A(_05652_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04517_)
  );
  OAI21X1 _11979_ (
    .A(_04298_),
    .B(_04505_),
    .C(_04517_),
    .Y(_04518_)
  );
  OAI21X1 _11980_ (
    .A( multiplier_0.reslo_3_ ),
    .B(_04507_),
    .C(_04518_),
    .Y(_04519_)
  );
  INVX1 _11981_ (
    .A(_04519_),
    .Y(_03968_)
  );
  AOI21X1 _11982_ (
    .A(_05653_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04520_)
  );
  OAI21X1 _11983_ (
    .A(_04308_),
    .B(_04505_),
    .C(_04520_),
    .Y(_04521_)
  );
  OAI21X1 _11984_ (
    .A( multiplier_0.reslo_4_ ),
    .B(_04507_),
    .C(_04521_),
    .Y(_04522_)
  );
  INVX1 _11985_ (
    .A(_04522_),
    .Y(_03969_)
  );
  AOI21X1 _11986_ (
    .A(_05654_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04523_)
  );
  OAI21X1 _11987_ (
    .A(_04318_),
    .B(_04505_),
    .C(_04523_),
    .Y(_04524_)
  );
  OAI21X1 _11988_ (
    .A( multiplier_0.reslo_5_ ),
    .B(_04507_),
    .C(_04524_),
    .Y(_04525_)
  );
  INVX1 _11989_ (
    .A(_04525_),
    .Y(_03970_)
  );
  AOI21X1 _11990_ (
    .A(_05655_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04526_)
  );
  OAI21X1 _11991_ (
    .A(_04327_),
    .B(_04505_),
    .C(_04526_),
    .Y(_04527_)
  );
  OAI21X1 _11992_ (
    .A( multiplier_0.reslo_6_ ),
    .B(_04507_),
    .C(_04527_),
    .Y(_04528_)
  );
  INVX1 _11993_ (
    .A(_04528_),
    .Y(_03971_)
  );
  AOI21X1 _11994_ (
    .A(_05656_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04529_)
  );
  OAI21X1 _11995_ (
    .A(_04337_),
    .B(_04505_),
    .C(_04529_),
    .Y(_04530_)
  );
  OAI21X1 _11996_ (
    .A( multiplier_0.reslo_7_ ),
    .B(_04507_),
    .C(_04530_),
    .Y(_04531_)
  );
  INVX1 _11997_ (
    .A(_04531_),
    .Y(_03972_)
  );
  AOI21X1 _11998_ (
    .A(_04464_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04532_)
  );
  OAI21X1 _11999_ (
    .A(_04346_),
    .B(_04505_),
    .C(_04532_),
    .Y(_04533_)
  );
  OAI21X1 _12000_ (
    .A( multiplier_0.reslo_8_ ),
    .B(_04507_),
    .C(_04533_),
    .Y(_04534_)
  );
  INVX1 _12001_ (
    .A(_04534_),
    .Y(_03973_)
  );
  AOI21X1 _12002_ (
    .A(_04469_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04535_)
  );
  OAI21X1 _12003_ (
    .A(_04356_),
    .B(_04505_),
    .C(_04535_),
    .Y(_04536_)
  );
  OAI21X1 _12004_ (
    .A( multiplier_0.reslo_9_ ),
    .B(_04507_),
    .C(_04536_),
    .Y(_04537_)
  );
  INVX1 _12005_ (
    .A(_04537_),
    .Y(_03974_)
  );
  AOI21X1 _12006_ (
    .A(_04474_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04538_)
  );
  OAI21X1 _12007_ (
    .A(_04365_),
    .B(_04505_),
    .C(_04538_),
    .Y(_04539_)
  );
  OAI21X1 _12008_ (
    .A( multiplier_0.reslo_10_ ),
    .B(_04507_),
    .C(_04539_),
    .Y(_04540_)
  );
  INVX1 _12009_ (
    .A(_04540_),
    .Y(_03975_)
  );
  AOI21X1 _12010_ (
    .A(_04479_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04541_)
  );
  OAI21X1 _12011_ (
    .A(_04374_),
    .B(_04505_),
    .C(_04541_),
    .Y(_04542_)
  );
  OAI21X1 _12012_ (
    .A( multiplier_0.reslo_11_ ),
    .B(_04507_),
    .C(_04542_),
    .Y(_04543_)
  );
  INVX1 _12013_ (
    .A(_04543_),
    .Y(_03976_)
  );
  AOI21X1 _12014_ (
    .A(_04484_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04544_)
  );
  OAI21X1 _12015_ (
    .A(_04383_),
    .B(_04505_),
    .C(_04544_),
    .Y(_04545_)
  );
  OAI21X1 _12016_ (
    .A( multiplier_0.reslo_12_ ),
    .B(_04507_),
    .C(_04545_),
    .Y(_04546_)
  );
  INVX1 _12017_ (
    .A(_04546_),
    .Y(_03977_)
  );
  AOI21X1 _12018_ (
    .A(_04489_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04547_)
  );
  OAI21X1 _12019_ (
    .A(_04393_),
    .B(_04505_),
    .C(_04547_),
    .Y(_04548_)
  );
  OAI21X1 _12020_ (
    .A( multiplier_0.reslo_13_ ),
    .B(_04507_),
    .C(_04548_),
    .Y(_04549_)
  );
  INVX1 _12021_ (
    .A(_04549_),
    .Y(_03978_)
  );
  AOI21X1 _12022_ (
    .A(_04494_),
    .B(_04503_),
    .C(_04506_),
    .Y(_04550_)
  );
  OAI21X1 _12023_ (
    .A(_04402_),
    .B(_04505_),
    .C(_04550_),
    .Y(_04551_)
  );
  OAI21X1 _12024_ (
    .A( multiplier_0.reslo_14_ ),
    .B(_04507_),
    .C(_04551_),
    .Y(_04552_)
  );
  INVX1 _12025_ (
    .A(_04552_),
    .Y(_03979_)
  );
  NOR2X1 _12026_ (
    .A(_04411_),
    .B(_04505_),
    .Y(_04553_)
  );
  OAI21X1 _12027_ (
    .A(_04499_),
    .B(_04504_),
    .C(_04507_),
    .Y(_04554_)
  );
  OAI22X1 _12028_ (
    .A( multiplier_0.reslo_15_ ),
    .B(_04507_),
    .C(_04553_),
    .D(_04554_),
    .Y(_04555_)
  );
  INVX1 _12029_ (
    .A(_04555_),
    .Y(_03980_)
  );
  MUX2X1 _12030_ (
    .A( multiplier_0.op2_0_ ),
    .B(_05643_),
    .S(_04429_),
    .Y(_04556_)
  );
  INVX1 _12031_ (
    .A(_04556_),
    .Y(_03981_)
  );
  MUX2X1 _12032_ (
    .A( multiplier_0.op2_1_ ),
    .B(_05650_),
    .S(_04429_),
    .Y(_04557_)
  );
  INVX1 _12033_ (
    .A(_04557_),
    .Y(_03982_)
  );
  MUX2X1 _12034_ (
    .A( multiplier_0.op2_2_ ),
    .B(_05651_),
    .S(_04429_),
    .Y(_04558_)
  );
  INVX1 _12035_ (
    .A(_04558_),
    .Y(_03983_)
  );
  MUX2X1 _12036_ (
    .A( multiplier_0.op2_3_ ),
    .B(_05652_),
    .S(_04429_),
    .Y(_04559_)
  );
  INVX1 _12037_ (
    .A(_04559_),
    .Y(_03984_)
  );
  MUX2X1 _12038_ (
    .A( multiplier_0.op2_4_ ),
    .B(_05653_),
    .S(_04429_),
    .Y(_04560_)
  );
  INVX1 _12039_ (
    .A(_04560_),
    .Y(_03985_)
  );
  MUX2X1 _12040_ (
    .A( multiplier_0.op2_5_ ),
    .B(_05654_),
    .S(_04429_),
    .Y(_04561_)
  );
  INVX1 _12041_ (
    .A(_04561_),
    .Y(_03986_)
  );
  MUX2X1 _12042_ (
    .A( multiplier_0.op2_6_ ),
    .B(_05655_),
    .S(_04429_),
    .Y(_04562_)
  );
  INVX1 _12043_ (
    .A(_04562_),
    .Y(_03987_)
  );
  MUX2X1 _12044_ (
    .A( multiplier_0.op2_7_ ),
    .B(_05656_),
    .S(_04429_),
    .Y(_04563_)
  );
  INVX1 _12045_ (
    .A(_04563_),
    .Y(_03988_)
  );
  OAI21X1 _12046_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_8_ ),
    .Y(_04564_)
  );
  OAI21X1 _12047_ (
    .A(_04429_),
    .B(_04465_),
    .C(_04564_),
    .Y(_03989_)
  );
  OAI21X1 _12048_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_9_ ),
    .Y(_04565_)
  );
  OAI21X1 _12049_ (
    .A(_04429_),
    .B(_04470_),
    .C(_04565_),
    .Y(_03990_)
  );
  OAI21X1 _12050_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_10_ ),
    .Y(_04566_)
  );
  OAI21X1 _12051_ (
    .A(_04429_),
    .B(_04475_),
    .C(_04566_),
    .Y(_03991_)
  );
  OAI21X1 _12052_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_11_ ),
    .Y(_04567_)
  );
  OAI21X1 _12053_ (
    .A(_04429_),
    .B(_04480_),
    .C(_04567_),
    .Y(_03992_)
  );
  OAI21X1 _12054_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_12_ ),
    .Y(_04568_)
  );
  OAI21X1 _12055_ (
    .A(_04429_),
    .B(_04485_),
    .C(_04568_),
    .Y(_03993_)
  );
  OAI21X1 _12056_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_13_ ),
    .Y(_04569_)
  );
  OAI21X1 _12057_ (
    .A(_04429_),
    .B(_04490_),
    .C(_04569_),
    .Y(_03994_)
  );
  OAI21X1 _12058_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_14_ ),
    .Y(_04570_)
  );
  OAI21X1 _12059_ (
    .A(_04429_),
    .B(_04495_),
    .C(_04570_),
    .Y(_03995_)
  );
  OAI21X1 _12060_ (
    .A(_04631_),
    .B(_04633_),
    .C( multiplier_0.op2_15_ ),
    .Y(_04571_)
  );
  OAI21X1 _12061_ (
    .A(_04429_),
    .B(_04499_),
    .C(_04571_),
    .Y(_03996_)
  );
  MUX2X1 _12062_ (
    .A( multiplier_0.op1_0_ ),
    .B(_05643_),
    .S(_04424_),
    .Y(_04572_)
  );
  INVX1 _12063_ (
    .A(_04572_),
    .Y(_03997_)
  );
  MUX2X1 _12064_ (
    .A( multiplier_0.op1_1_ ),
    .B(_05650_),
    .S(_04424_),
    .Y(_04573_)
  );
  INVX1 _12065_ (
    .A(_04573_),
    .Y(_03998_)
  );
  MUX2X1 _12066_ (
    .A( multiplier_0.op1_2_ ),
    .B(_05651_),
    .S(_04424_),
    .Y(_04574_)
  );
  INVX1 _12067_ (
    .A(_04574_),
    .Y(_03999_)
  );
  MUX2X1 _12068_ (
    .A( multiplier_0.op1_3_ ),
    .B(_05652_),
    .S(_04424_),
    .Y(_04575_)
  );
  INVX1 _12069_ (
    .A(_04575_),
    .Y(_04000_)
  );
  MUX2X1 _12070_ (
    .A( multiplier_0.op1_4_ ),
    .B(_05653_),
    .S(_04424_),
    .Y(_04576_)
  );
  INVX1 _12071_ (
    .A(_04576_),
    .Y(_04001_)
  );
  MUX2X1 _12072_ (
    .A( multiplier_0.op1_5_ ),
    .B(_05654_),
    .S(_04424_),
    .Y(_04577_)
  );
  INVX1 _12073_ (
    .A(_04577_),
    .Y(_04002_)
  );
  MUX2X1 _12074_ (
    .A( multiplier_0.op1_6_ ),
    .B(_05655_),
    .S(_04424_),
    .Y(_04578_)
  );
  INVX1 _12075_ (
    .A(_04578_),
    .Y(_04003_)
  );
  MUX2X1 _12076_ (
    .A( multiplier_0.op1_7_ ),
    .B(_05656_),
    .S(_04424_),
    .Y(_04579_)
  );
  INVX1 _12077_ (
    .A(_04579_),
    .Y(_04004_)
  );
  OAI21X1 _12078_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_8_ ),
    .Y(_04580_)
  );
  OAI21X1 _12079_ (
    .A(_04424_),
    .B(_04465_),
    .C(_04580_),
    .Y(_04005_)
  );
  OAI21X1 _12080_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_9_ ),
    .Y(_04581_)
  );
  OAI21X1 _12081_ (
    .A(_04424_),
    .B(_04470_),
    .C(_04581_),
    .Y(_04006_)
  );
  OAI21X1 _12082_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_10_ ),
    .Y(_04582_)
  );
  OAI21X1 _12083_ (
    .A(_04424_),
    .B(_04475_),
    .C(_04582_),
    .Y(_04007_)
  );
  OAI21X1 _12084_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_11_ ),
    .Y(_04583_)
  );
  OAI21X1 _12085_ (
    .A(_04424_),
    .B(_04480_),
    .C(_04583_),
    .Y(_04008_)
  );
  OAI21X1 _12086_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_12_ ),
    .Y(_04584_)
  );
  OAI21X1 _12087_ (
    .A(_04424_),
    .B(_04485_),
    .C(_04584_),
    .Y(_04009_)
  );
  OAI21X1 _12088_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_13_ ),
    .Y(_04585_)
  );
  OAI21X1 _12089_ (
    .A(_04424_),
    .B(_04490_),
    .C(_04585_),
    .Y(_04010_)
  );
  OAI21X1 _12090_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_14_ ),
    .Y(_04586_)
  );
  OAI21X1 _12091_ (
    .A(_04424_),
    .B(_04495_),
    .C(_04586_),
    .Y(_04011_)
  );
  OAI21X1 _12092_ (
    .A(_05635_),
    .B(_04631_),
    .C( multiplier_0.op1_15_ ),
    .Y(_04587_)
  );
  OAI21X1 _12093_ (
    .A(_04424_),
    .B(_04499_),
    .C(_04587_),
    .Y(_04012_)
  );
  DFFSR _12094_ (
    .CLK(dco_clk),
    .D( multiplier_0.op2_wr ),
    .Q( multiplier_0.cycle_0_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12095_ (
    .CLK(dco_clk),
    .D( multiplier_0.cycle_0_ ),
    .Q( multiplier_0.cycle_1_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12096_ (
    .CLK(dco_clk),
    .D(_03945_),
    .Q( multiplier_0.acc_sel ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12097_ (
    .CLK(dco_clk),
    .D(_03946_),
    .Q( multiplier_0.sign_sel ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12098_ (
    .CLK(dco_clk),
    .D(_03947_),
    .Q( multiplier_0.sumext_0_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12099_ (
    .CLK(dco_clk),
    .D(_03948_),
    .Q( multiplier_0.sumext_10_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12100_ (
    .CLK(dco_clk),
    .D(_03949_),
    .Q( multiplier_0.reshi_0_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12101_ (
    .CLK(dco_clk),
    .D(_03950_),
    .Q( multiplier_0.reshi_1_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12102_ (
    .CLK(dco_clk),
    .D(_03951_),
    .Q( multiplier_0.reshi_2_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12103_ (
    .CLK(dco_clk),
    .D(_03952_),
    .Q( multiplier_0.reshi_3_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12104_ (
    .CLK(dco_clk),
    .D(_03953_),
    .Q( multiplier_0.reshi_4_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12105_ (
    .CLK(dco_clk),
    .D(_03954_),
    .Q( multiplier_0.reshi_5_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12106_ (
    .CLK(dco_clk),
    .D(_03955_),
    .Q( multiplier_0.reshi_6_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12107_ (
    .CLK(dco_clk),
    .D(_03956_),
    .Q( multiplier_0.reshi_7_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12108_ (
    .CLK(dco_clk),
    .D(_03957_),
    .Q( multiplier_0.reshi_8_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12109_ (
    .CLK(dco_clk),
    .D(_03958_),
    .Q( multiplier_0.reshi_9_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12110_ (
    .CLK(dco_clk),
    .D(_03959_),
    .Q( multiplier_0.reshi_10_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12111_ (
    .CLK(dco_clk),
    .D(_03960_),
    .Q( multiplier_0.reshi_11_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12112_ (
    .CLK(dco_clk),
    .D(_03961_),
    .Q( multiplier_0.reshi_12_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12113_ (
    .CLK(dco_clk),
    .D(_03962_),
    .Q( multiplier_0.reshi_13_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12114_ (
    .CLK(dco_clk),
    .D(_03963_),
    .Q( multiplier_0.reshi_14_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12115_ (
    .CLK(dco_clk),
    .D(_03964_),
    .Q( multiplier_0.reshi_15_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12116_ (
    .CLK(dco_clk),
    .D(_03965_),
    .Q( multiplier_0.reslo_0_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12117_ (
    .CLK(dco_clk),
    .D(_03966_),
    .Q( multiplier_0.reslo_1_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12118_ (
    .CLK(dco_clk),
    .D(_03967_),
    .Q( multiplier_0.reslo_2_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12119_ (
    .CLK(dco_clk),
    .D(_03968_),
    .Q( multiplier_0.reslo_3_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12120_ (
    .CLK(dco_clk),
    .D(_03969_),
    .Q( multiplier_0.reslo_4_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12121_ (
    .CLK(dco_clk),
    .D(_03970_),
    .Q( multiplier_0.reslo_5_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12122_ (
    .CLK(dco_clk),
    .D(_03971_),
    .Q( multiplier_0.reslo_6_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12123_ (
    .CLK(dco_clk),
    .D(_03972_),
    .Q( multiplier_0.reslo_7_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12124_ (
    .CLK(dco_clk),
    .D(_03973_),
    .Q( multiplier_0.reslo_8_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12125_ (
    .CLK(dco_clk),
    .D(_03974_),
    .Q( multiplier_0.reslo_9_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12126_ (
    .CLK(dco_clk),
    .D(_03975_),
    .Q( multiplier_0.reslo_10_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12127_ (
    .CLK(dco_clk),
    .D(_03976_),
    .Q( multiplier_0.reslo_11_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12128_ (
    .CLK(dco_clk),
    .D(_03977_),
    .Q( multiplier_0.reslo_12_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12129_ (
    .CLK(dco_clk),
    .D(_03978_),
    .Q( multiplier_0.reslo_13_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12130_ (
    .CLK(dco_clk),
    .D(_03979_),
    .Q( multiplier_0.reslo_14_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12131_ (
    .CLK(dco_clk),
    .D(_03980_),
    .Q( multiplier_0.reslo_15_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12132_ (
    .CLK(dco_clk),
    .D(_03981_),
    .Q( multiplier_0.op2_0_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12133_ (
    .CLK(dco_clk),
    .D(_03982_),
    .Q( multiplier_0.op2_1_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12134_ (
    .CLK(dco_clk),
    .D(_03983_),
    .Q( multiplier_0.op2_2_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12135_ (
    .CLK(dco_clk),
    .D(_03984_),
    .Q( multiplier_0.op2_3_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12136_ (
    .CLK(dco_clk),
    .D(_03985_),
    .Q( multiplier_0.op2_4_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12137_ (
    .CLK(dco_clk),
    .D(_03986_),
    .Q( multiplier_0.op2_5_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12138_ (
    .CLK(dco_clk),
    .D(_03987_),
    .Q( multiplier_0.op2_6_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12139_ (
    .CLK(dco_clk),
    .D(_03988_),
    .Q( multiplier_0.op2_7_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12140_ (
    .CLK(dco_clk),
    .D(_03989_),
    .Q( multiplier_0.op2_8_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12141_ (
    .CLK(dco_clk),
    .D(_03990_),
    .Q( multiplier_0.op2_9_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12142_ (
    .CLK(dco_clk),
    .D(_03991_),
    .Q( multiplier_0.op2_10_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12143_ (
    .CLK(dco_clk),
    .D(_03992_),
    .Q( multiplier_0.op2_11_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12144_ (
    .CLK(dco_clk),
    .D(_03993_),
    .Q( multiplier_0.op2_12_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12145_ (
    .CLK(dco_clk),
    .D(_03994_),
    .Q( multiplier_0.op2_13_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12146_ (
    .CLK(dco_clk),
    .D(_03995_),
    .Q( multiplier_0.op2_14_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12147_ (
    .CLK(dco_clk),
    .D(_03996_),
    .Q( multiplier_0.op2_15_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12148_ (
    .CLK(dco_clk),
    .D(_03997_),
    .Q( multiplier_0.op1_0_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12149_ (
    .CLK(dco_clk),
    .D(_03998_),
    .Q( multiplier_0.op1_1_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12150_ (
    .CLK(dco_clk),
    .D(_03999_),
    .Q( multiplier_0.op1_2_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12151_ (
    .CLK(dco_clk),
    .D(_04000_),
    .Q( multiplier_0.op1_3_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12152_ (
    .CLK(dco_clk),
    .D(_04001_),
    .Q( multiplier_0.op1_4_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12153_ (
    .CLK(dco_clk),
    .D(_04002_),
    .Q( multiplier_0.op1_5_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12154_ (
    .CLK(dco_clk),
    .D(_04003_),
    .Q( multiplier_0.op1_6_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12155_ (
    .CLK(dco_clk),
    .D(_04004_),
    .Q( multiplier_0.op1_7_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12156_ (
    .CLK(dco_clk),
    .D(_04005_),
    .Q( multiplier_0.op1_8_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12157_ (
    .CLK(dco_clk),
    .D(_04006_),
    .Q( multiplier_0.op1_9_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12158_ (
    .CLK(dco_clk),
    .D(_04007_),
    .Q( multiplier_0.op1_10_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12159_ (
    .CLK(dco_clk),
    .D(_04008_),
    .Q( multiplier_0.op1_11_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12160_ (
    .CLK(dco_clk),
    .D(_04009_),
    .Q( multiplier_0.op1_12_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12161_ (
    .CLK(dco_clk),
    .D(_04010_),
    .Q( multiplier_0.op1_13_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12162_ (
    .CLK(dco_clk),
    .D(_04011_),
    .Q( multiplier_0.op1_14_ ),
    .R(_03944_),
    .S(1'h1)
  );
  DFFSR _12163_ (
    .CLK(dco_clk),
    .D(_04012_),
    .Q( multiplier_0.op1_15_ ),
    .R(_03944_),
    .S(1'h1)
  );
  INVX1 _12164_ (
    .A(_05635_),
    .Y(_05403_)
  );
  INVX1 _12165_ (
    .A(_05633_),
    .Y(_05404_)
  );
  INVX1 _12166_ (
    .A(1'h0),
    .Y(_05405_)
  );
  INVX1 _12167_ (
    .A(1'h0),
    .Y(_05406_)
  );
  INVX1 _12168_ (
    .A(1'h0),
    .Y(_05407_)
  );
  INVX1 _12169_ (
    .A(1'h0),
    .Y(_05408_)
  );
  INVX1 _12170_ (
    .A( sfr_0.ie1_0_ ),
    .Y(_05409_)
  );
  INVX1 _12171_ (
    .A(_05643_),
    .Y(_05410_)
  );
  INVX1 _12172_ (
    .A(1'h0),
    .Y(_05411_)
  );
  INVX1 _12173_ (
    .A(1'h0),
    .Y(_05412_)
  );
  INVX1 _12174_ (
    .A(1'h0),
    .Y(_05413_)
  );
  INVX1 _12175_ (
    .A(1'h0),
    .Y(_05414_)
  );
  INVX1 _12176_ (
    .A(1'h0),
    .Y(_05415_)
  );
  INVX1 _12177_ (
    .A(1'h0),
    .Y(_05416_)
  );
  INVX1 _12178_ (
    .A(1'h0),
    .Y(_05417_)
  );
  INVX1 _12179_ (
    .A(1'h0),
    .Y(_05418_)
  );
  INVX1 _12180_ (
    .A(1'h0),
    .Y(_05419_)
  );
  INVX1 _12181_ (
    .A(1'h0),
    .Y(_05420_)
  );
  INVX1 _12182_ (
    .A(1'h0),
    .Y(_05421_)
  );
  INVX1 _12183_ (
    .A(_05695_),
    .Y(_05395_)
  );
  NOR2X1 _12184_ (
    .A(_05632_),
    .B(1'h0),
    .Y(_05422_)
  );
  NAND3X1 _12185_ (
    .A(_05404_),
    .B(_05659_),
    .C(_05422_),
    .Y(_05423_)
  );
  NOR2X1 _12186_ (
    .A(_05641_),
    .B(_05640_),
    .Y(_05424_)
  );
  NOR2X1 _12187_ (
    .A(_05631_),
    .B(_05642_),
    .Y(_05425_)
  );
  NAND2X1 _12188_ (
    .A(_05424_),
    .B(_05425_),
    .Y(_05426_)
  );
  NOR2X1 _12189_ (
    .A(_05637_),
    .B(_05636_),
    .Y(_05427_)
  );
  NOR2X1 _12190_ (
    .A(_05639_),
    .B(_05638_),
    .Y(_05428_)
  );
  NAND2X1 _12191_ (
    .A(_05427_),
    .B(_05428_),
    .Y(_05429_)
  );
  NOR3X1 _12192_ (
    .A(_05423_),
    .B(_05426_),
    .C(_05429_),
    .Y(_05430_)
  );
  NOR2X1 _12193_ (
    .A(_05661_),
    .B(_05660_),
    .Y(_05431_)
  );
  NAND2X1 _12194_ (
    .A(_05430_),
    .B(_05431_),
    .Y(_05432_)
  );
  NOR2X1 _12195_ (
    .A(_05630_),
    .B(_05634_),
    .Y(_05433_)
  );
  AND2X1 _12196_ (
    .A(_05635_),
    .B(_05433_),
    .Y(_05434_)
  );
  NAND3X1 _12197_ (
    .A(_05430_),
    .B(_05431_),
    .C(_05434_),
    .Y(_05435_)
  );
  NAND2X1 _12198_ (
    .A(_05403_),
    .B(_05634_),
    .Y(_05436_)
  );
  NOR2X1 _12199_ (
    .A(_05630_),
    .B(_05436_),
    .Y(_05437_)
  );
  NAND3X1 _12200_ (
    .A(_05430_),
    .B(_05431_),
    .C(_05437_),
    .Y(_05438_)
  );
  OAI21X1 _12201_ (
    .A(_05405_),
    .B(_05435_),
    .C(_05438_),
    .Y( sfr_0.per_dout_14_ )
  );
  NAND2X1 _12202_ (
    .A(_05403_),
    .B(_05630_),
    .Y(_05439_)
  );
  NAND3X1 _12203_ (
    .A(_05403_),
    .B(_05630_),
    .C(_05634_),
    .Y(_05440_)
  );
  INVX1 _12204_ (
    .A(_05440_),
    .Y(_05441_)
  );
  NAND3X1 _12205_ (
    .A(_05430_),
    .B(_05431_),
    .C(_05441_),
    .Y(_05442_)
  );
  OAI21X1 _12206_ (
    .A(_05406_),
    .B(_05435_),
    .C(_05442_),
    .Y( sfr_0.per_dout_8_ )
  );
  OAI21X1 _12207_ (
    .A(_05407_),
    .B(_05435_),
    .C(_05442_),
    .Y( sfr_0.per_dout_15_ )
  );
  OAI21X1 _12208_ (
    .A(_05408_),
    .B(_05435_),
    .C(_05438_),
    .Y( sfr_0.per_dout_1_ )
  );
  AND2X1 _12209_ (
    .A(_05403_),
    .B(_05433_),
    .Y(_05397_)
  );
  AOI22X1 _12210_ (
    .A(_05403_),
    .B(_05634_),
    .C( sfr_0.ie1_0_ ),
    .D(_05397_),
    .Y(_05398_)
  );
  NOR2X1 _12211_ (
    .A(_05634_),
    .B(_05439_),
    .Y(_05399_)
  );
  AOI22X1 _12212_ (
    .A(1'h0),
    .B(_05434_),
    .C(_05399_),
    .D( sfr_0.ifg1_0_ ),
    .Y(_05400_)
  );
  AOI21X1 _12213_ (
    .A(_05398_),
    .B(_05400_),
    .C(_05432_),
    .Y( sfr_0.per_dout_0_ )
  );
  NAND3X1 _12214_ (
    .A(_05660_),
    .B(_05430_),
    .C(_05399_),
    .Y(_05401_)
  );
  NOR2X1 _12215_ (
    .A(_05643_),
    .B(_05401_),
    .Y( sfr_0.wdtifg_sw_clr )
  );
  NOR2X1 _12216_ (
    .A(_05410_),
    .B(_05401_),
    .Y( sfr_0.wdtifg_sw_set )
  );
  NOR2X1 _12217_ (
    .A(_05411_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_2_ )
  );
  NOR2X1 _12218_ (
    .A(_05412_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_3_ )
  );
  NOR2X1 _12219_ (
    .A(_05413_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_4_ )
  );
  NOR2X1 _12220_ (
    .A(_05414_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_5_ )
  );
  NOR2X1 _12221_ (
    .A(_05415_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_6_ )
  );
  NOR2X1 _12222_ (
    .A(_05416_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_7_ )
  );
  NOR2X1 _12223_ (
    .A(_05417_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_9_ )
  );
  NOR2X1 _12224_ (
    .A(_05418_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_10_ )
  );
  NOR2X1 _12225_ (
    .A(_05419_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_11_ )
  );
  NOR2X1 _12226_ (
    .A(_05420_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_12_ )
  );
  NOR2X1 _12227_ (
    .A(_05421_),
    .B(_05435_),
    .Y( sfr_0.cpu_nr_rd_13_ )
  );
  NAND3X1 _12228_ (
    .A(_05660_),
    .B(_05430_),
    .C(_05397_),
    .Y(_05402_)
  );
  MUX2X1 _12229_ (
    .A(_05409_),
    .B(_05410_),
    .S(_05402_),
    .Y(_05396_)
  );
  DFFSR _12230_ (
    .CLK(dco_clk),
    .D(_05396_),
    .Q( sfr_0.ie1_0_ ),
    .R(_05395_),
    .S(1'h1)
  );
  INVX1 _12231_ (
    .A( watchdog_0.wdtcnt_2_ ),
    .Y(_05576_)
  );
  INVX1 _12232_ (
    .A( watchdog_0.wdtctl_0_ ),
    .Y(_05577_)
  );
  INVX1 _12233_ (
    .A( watchdog_0.wdtctl_1_ ),
    .Y(_05578_)
  );
  INVX1 _12234_ (
    .A( watchdog_0.wdtcnt_9_ ),
    .Y(_05579_)
  );
  INVX1 _12235_ (
    .A( watchdog_0.wdtcnt_10_ ),
    .Y(_05580_)
  );
  INVX1 _12236_ (
    .A(_05639_),
    .Y(_05468_)
  );
  INVX1 _12237_ (
    .A(_05641_),
    .Y(_05469_)
  );
  INVX1 _12238_ (
    .A(_05631_),
    .Y(_05470_)
  );
  INVX1 _12239_ (
    .A(_05633_),
    .Y(_05471_)
  );
  INVX1 _12240_ (
    .A(_05659_),
    .Y(_05472_)
  );
  INVX1 _12241_ (
    .A( sfr_0.wdtifg_sw_set ),
    .Y(_05473_)
  );
  INVX1 _12242_ (
    .A( sfr_0.wdtifg_sw_clr ),
    .Y(_05474_)
  );
  INVX1 _12243_ (
    .A( clock_module_0.por ),
    .Y(_05444_)
  );
  INVX1 _12244_ (
    .A(_05695_),
    .Y(_05445_)
  );
  NOR2X1 _12245_ (
    .A(_05661_),
    .B(_05660_),
    .Y(_05475_)
  );
  NOR2X1 _12246_ (
    .A(_05638_),
    .B(_05641_),
    .Y(_05476_)
  );
  NAND3X1 _12247_ (
    .A(_05637_),
    .B(_05468_),
    .C(_05476_),
    .Y(_05477_)
  );
  NOR2X1 _12248_ (
    .A(_05630_),
    .B(_05635_),
    .Y(_05478_)
  );
  NOR2X1 _12249_ (
    .A(_05634_),
    .B(_05636_),
    .Y(_05479_)
  );
  NAND2X1 _12250_ (
    .A(_05478_),
    .B(_05479_),
    .Y(_05480_)
  );
  NOR2X1 _12251_ (
    .A(_05477_),
    .B(_05480_),
    .Y(_05481_)
  );
  NOR2X1 _12252_ (
    .A(_05632_),
    .B(1'h0),
    .Y(_05482_)
  );
  NAND2X1 _12253_ (
    .A(_05659_),
    .B(_05482_),
    .Y(_05483_)
  );
  NOR2X1 _12254_ (
    .A(_05642_),
    .B(_05633_),
    .Y(_05484_)
  );
  NAND3X1 _12255_ (
    .A(_05640_),
    .B(_05470_),
    .C(_05484_),
    .Y(_05485_)
  );
  NOR2X1 _12256_ (
    .A(_05483_),
    .B(_05485_),
    .Y(_05486_)
  );
  NAND3X1 _12257_ (
    .A(_05475_),
    .B(_05481_),
    .C(_05486_),
    .Y(_05487_)
  );
  INVX1 _12258_ (
    .A(_05487_),
    .Y( watchdog_0.per_dout_11_ )
  );
  NOR2X1 _12259_ (
    .A(_05577_),
    .B(_05487_),
    .Y( watchdog_0.per_dout_0_ )
  );
  NOR2X1 _12260_ (
    .A(_05578_),
    .B(_05487_),
    .Y( watchdog_0.per_dout_1_ )
  );
  AND2X1 _12261_ (
    .A( watchdog_0.wdtctl_2_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_2_ )
  );
  AND2X1 _12262_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_4_ )
  );
  AND2X1 _12263_ (
    .A( watchdog_0.wdtctl_7_ ),
    .B( watchdog_0.per_dout_11_ ),
    .Y( watchdog_0.per_dout_7_ )
  );
  NAND3X1 _12264_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B( sfr_0.ifg1_0_ ),
    .C( sfr_0.ie1_0_ ),
    .Y(_05488_)
  );
  INVX1 _12265_ (
    .A(_05488_),
    .Y( frontend_0.wdt_irq )
  );
  MUX2X1 _12266_ (
    .A(_05581_),
    .B(_05696_),
    .S( watchdog_0.wdtctl_2_ ),
    .Y(_05489_)
  );
  OR2X1 _12267_ (
    .A( watchdog_0.wdtctl_7_ ),
    .B(_05582_),
    .Y(_05490_)
  );
  NOR2X1 _12268_ (
    .A(_05489_),
    .B(_05490_),
    .Y(_05491_)
  );
  INVX1 _12269_ (
    .A(_05491_),
    .Y(_05492_)
  );
  NOR2X1 _12270_ (
    .A( watchdog_0.wdtctl_0_ ),
    .B( watchdog_0.wdtctl_1_ ),
    .Y(_05493_)
  );
  NAND2X1 _12271_ (
    .A( watchdog_0.wdtcnt_5_ ),
    .B( watchdog_0.wdtcnt_4_ ),
    .Y(_05494_)
  );
  NAND2X1 _12272_ (
    .A( watchdog_0.wdtcnt_1_ ),
    .B( watchdog_0.wdtcnt_0_ ),
    .Y(_05495_)
  );
  NAND2X1 _12273_ (
    .A( watchdog_0.wdtcnt_3_ ),
    .B( watchdog_0.wdtcnt_2_ ),
    .Y(_05496_)
  );
  NOR3X1 _12274_ (
    .A(_05494_),
    .B(_05495_),
    .C(_05496_),
    .Y(_05497_)
  );
  AND2X1 _12275_ (
    .A( watchdog_0.wdtcnt_7_ ),
    .B( watchdog_0.wdtcnt_8_ ),
    .Y(_05498_)
  );
  NAND3X1 _12276_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B(_05497_),
    .C(_05498_),
    .Y(_05499_)
  );
  NOR2X1 _12277_ (
    .A(_05579_),
    .B(_05499_),
    .Y(_05500_)
  );
  XNOR2X1 _12278_ (
    .A(_05579_),
    .B(_05499_),
    .Y(_05501_)
  );
  NAND3X1 _12279_ (
    .A( watchdog_0.wdtcnt_11_ ),
    .B( watchdog_0.wdtcnt_10_ ),
    .C( watchdog_0.wdtcnt_12_ ),
    .Y(_05502_)
  );
  NOR3X1 _12280_ (
    .A(_05579_),
    .B(_05499_),
    .C(_05502_),
    .Y(_05503_)
  );
  XOR2X1 _12281_ (
    .A( watchdog_0.wdtcnt_13_ ),
    .B(_05503_),
    .Y(_05504_)
  );
  OAI21X1 _12282_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B(_05497_),
    .C( watchdog_0.wdtctl_1_ ),
    .Y(_05505_)
  );
  OR2X1 _12283_ (
    .A(_05577_),
    .B(_05505_),
    .Y(_05506_)
  );
  AOI21X1 _12284_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B(_05497_),
    .C(_05506_),
    .Y(_05507_)
  );
  NAND3X1 _12285_ (
    .A( watchdog_0.wdtcnt_13_ ),
    .B( watchdog_0.wdtcnt_14_ ),
    .C(_05503_),
    .Y(_05508_)
  );
  XOR2X1 _12286_ (
    .A( watchdog_0.wdtcnt_15_ ),
    .B(_05508_),
    .Y(_05509_)
  );
  AOI21X1 _12287_ (
    .A( watchdog_0.wdtctl_1_ ),
    .B(_05501_),
    .C( watchdog_0.wdtctl_0_ ),
    .Y(_05510_)
  );
  AOI21X1 _12288_ (
    .A(_05578_),
    .B(_05504_),
    .C(_05510_),
    .Y(_05511_)
  );
  AOI21X1 _12289_ (
    .A(_05493_),
    .B(_05509_),
    .C(_05511_),
    .Y(_05512_)
  );
  OAI21X1 _12290_ (
    .A(_05507_),
    .B(_05512_),
    .C(_05491_),
    .Y(_05513_)
  );
  NOR2X1 _12291_ (
    .A(_05639_),
    .B(_05638_),
    .Y(_05514_)
  );
  NOR2X1 _12292_ (
    .A(_05630_),
    .B(_05636_),
    .Y(_05515_)
  );
  OR2X1 _12293_ (
    .A(_05631_),
    .B(_05642_),
    .Y(_05516_)
  );
  NOR2X1 _12294_ (
    .A(_05632_),
    .B(_05516_),
    .Y(_05517_)
  );
  NAND3X1 _12295_ (
    .A(_05514_),
    .B(_05515_),
    .C(_05517_),
    .Y(_05518_)
  );
  NOR2X1 _12296_ (
    .A(_05635_),
    .B(_05634_),
    .Y(_05519_)
  );
  NAND3X1 _12297_ (
    .A(_05637_),
    .B(_05469_),
    .C(_05519_),
    .Y(_05520_)
  );
  NOR2X1 _12298_ (
    .A(1'h0),
    .B(_05472_),
    .Y(_05521_)
  );
  NAND3X1 _12299_ (
    .A(_05640_),
    .B(_05471_),
    .C(_05521_),
    .Y(_05522_)
  );
  OR2X1 _12300_ (
    .A(_05520_),
    .B(_05522_),
    .Y(_05523_)
  );
  NOR2X1 _12301_ (
    .A(_05518_),
    .B(_05523_),
    .Y(_05524_)
  );
  OAI21X1 _12302_ (
    .A(_05661_),
    .B(_05660_),
    .C(_05524_),
    .Y(_05525_)
  );
  INVX1 _12303_ (
    .A(_05525_),
    .Y(_05526_)
  );
  OR2X1 _12304_ (
    .A(_05647_),
    .B(_05649_),
    .Y(_05527_)
  );
  NOR2X1 _12305_ (
    .A(_05657_),
    .B(_05644_),
    .Y(_05528_)
  );
  NAND3X1 _12306_ (
    .A(_05646_),
    .B(_05648_),
    .C(_05528_),
    .Y(_05529_)
  );
  INVX1 _12307_ (
    .A(_05529_),
    .Y(_05530_)
  );
  NAND3X1 _12308_ (
    .A(_05658_),
    .B(_05645_),
    .C(_05530_),
    .Y(_05531_)
  );
  OAI21X1 _12309_ (
    .A(_05527_),
    .B(_05531_),
    .C(_05526_),
    .Y(_05532_)
  );
  AND2X1 _12310_ (
    .A(_05513_),
    .B(_05532_),
    .Y(_05533_)
  );
  AOI22X1 _12311_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B(_05532_),
    .C(_05533_),
    .D(_05473_),
    .Y(_05443_)
  );
  MUX2X1 _12312_ (
    .A( watchdog_0.wdtctl_0_ ),
    .B(_05643_),
    .S(_05525_),
    .Y(_05534_)
  );
  INVX1 _12313_ (
    .A(_05534_),
    .Y(_05446_)
  );
  MUX2X1 _12314_ (
    .A( watchdog_0.wdtctl_1_ ),
    .B(_05650_),
    .S(_05525_),
    .Y(_05535_)
  );
  INVX1 _12315_ (
    .A(_05535_),
    .Y(_05447_)
  );
  MUX2X1 _12316_ (
    .A( watchdog_0.wdtctl_2_ ),
    .B(_05651_),
    .S(_05525_),
    .Y(_05536_)
  );
  INVX1 _12317_ (
    .A(_05536_),
    .Y(_05448_)
  );
  MUX2X1 _12318_ (
    .A( watchdog_0.wdtctl_4_ ),
    .B(_05653_),
    .S(_05525_),
    .Y(_05537_)
  );
  INVX1 _12319_ (
    .A(_05537_),
    .Y(_05449_)
  );
  MUX2X1 _12320_ (
    .A( watchdog_0.wdtctl_7_ ),
    .B(_05656_),
    .S(_05525_),
    .Y(_05538_)
  );
  INVX1 _12321_ (
    .A(_05538_),
    .Y(_05450_)
  );
  NAND2X1 _12322_ (
    .A(_05617_),
    .B( watchdog_0.wdtctl_4_ ),
    .Y(_05539_)
  );
  NAND3X1 _12323_ (
    .A(_05474_),
    .B( sfr_0.ifg1_0_ ),
    .C(_05539_),
    .Y(_05540_)
  );
  NAND3X1 _12324_ (
    .A(_05473_),
    .B(_05533_),
    .C(_05540_),
    .Y(_05451_)
  );
  NAND2X1 _12325_ (
    .A(_05652_),
    .B(_05526_),
    .Y(_05541_)
  );
  NAND3X1 _12326_ (
    .A(_05513_),
    .B(_05532_),
    .C(_05541_),
    .Y(_05542_)
  );
  NAND2X1 _12327_ (
    .A( watchdog_0.wdtcnt_0_ ),
    .B(_05491_),
    .Y(_05543_)
  );
  XNOR2X1 _12328_ (
    .A( watchdog_0.wdtcnt_0_ ),
    .B(_05491_),
    .Y(_05544_)
  );
  NOR2X1 _12329_ (
    .A(_05542_),
    .B(_05544_),
    .Y(_05452_)
  );
  OR2X1 _12330_ (
    .A(_05492_),
    .B(_05495_),
    .Y(_05545_)
  );
  XOR2X1 _12331_ (
    .A( watchdog_0.wdtcnt_1_ ),
    .B(_05543_),
    .Y(_05546_)
  );
  NOR2X1 _12332_ (
    .A(_05542_),
    .B(_05546_),
    .Y(_05453_)
  );
  NOR2X1 _12333_ (
    .A(_05576_),
    .B(_05545_),
    .Y(_05547_)
  );
  XNOR2X1 _12334_ (
    .A(_05576_),
    .B(_05545_),
    .Y(_05548_)
  );
  NOR2X1 _12335_ (
    .A(_05542_),
    .B(_05548_),
    .Y(_05454_)
  );
  XNOR2X1 _12336_ (
    .A( watchdog_0.wdtcnt_3_ ),
    .B(_05547_),
    .Y(_05549_)
  );
  NOR2X1 _12337_ (
    .A(_05542_),
    .B(_05549_),
    .Y(_05455_)
  );
  AOI21X1 _12338_ (
    .A( watchdog_0.wdtcnt_3_ ),
    .B(_05547_),
    .C( watchdog_0.wdtcnt_4_ ),
    .Y(_05550_)
  );
  NAND3X1 _12339_ (
    .A( watchdog_0.wdtcnt_4_ ),
    .B( watchdog_0.wdtcnt_3_ ),
    .C(_05547_),
    .Y(_05551_)
  );
  INVX1 _12340_ (
    .A(_05551_),
    .Y(_05552_)
  );
  NOR3X1 _12341_ (
    .A(_05542_),
    .B(_05550_),
    .C(_05552_),
    .Y(_05456_)
  );
  AND2X1 _12342_ (
    .A(_05491_),
    .B(_05497_),
    .Y(_05553_)
  );
  INVX1 _12343_ (
    .A(_05553_),
    .Y(_05554_)
  );
  OAI21X1 _12344_ (
    .A( watchdog_0.wdtcnt_5_ ),
    .B(_05552_),
    .C(_05554_),
    .Y(_05555_)
  );
  NOR2X1 _12345_ (
    .A(_05542_),
    .B(_05555_),
    .Y(_05457_)
  );
  NAND2X1 _12346_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B(_05553_),
    .Y(_05556_)
  );
  XNOR2X1 _12347_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B(_05553_),
    .Y(_05557_)
  );
  NOR2X1 _12348_ (
    .A(_05542_),
    .B(_05557_),
    .Y(_05458_)
  );
  NAND3X1 _12349_ (
    .A( watchdog_0.wdtcnt_6_ ),
    .B( watchdog_0.wdtcnt_7_ ),
    .C(_05553_),
    .Y(_05558_)
  );
  XOR2X1 _12350_ (
    .A( watchdog_0.wdtcnt_7_ ),
    .B(_05556_),
    .Y(_05559_)
  );
  NOR2X1 _12351_ (
    .A(_05542_),
    .B(_05559_),
    .Y(_05459_)
  );
  XOR2X1 _12352_ (
    .A( watchdog_0.wdtcnt_8_ ),
    .B(_05558_),
    .Y(_05560_)
  );
  NOR2X1 _12353_ (
    .A(_05542_),
    .B(_05560_),
    .Y(_05460_)
  );
  NAND2X1 _12354_ (
    .A(_05491_),
    .B(_05501_),
    .Y(_05561_)
  );
  OAI21X1 _12355_ (
    .A( watchdog_0.wdtcnt_9_ ),
    .B(_05491_),
    .C(_05561_),
    .Y(_05562_)
  );
  NOR2X1 _12356_ (
    .A(_05542_),
    .B(_05562_),
    .Y(_05461_)
  );
  NAND2X1 _12357_ (
    .A(_05491_),
    .B(_05500_),
    .Y(_05563_)
  );
  AOI21X1 _12358_ (
    .A(_05491_),
    .B(_05500_),
    .C( watchdog_0.wdtcnt_10_ ),
    .Y(_05564_)
  );
  NOR2X1 _12359_ (
    .A(_05580_),
    .B(_05563_),
    .Y(_05565_)
  );
  NOR3X1 _12360_ (
    .A(_05542_),
    .B(_05564_),
    .C(_05565_),
    .Y(_05462_)
  );
  XNOR2X1 _12361_ (
    .A( watchdog_0.wdtcnt_11_ ),
    .B(_05565_),
    .Y(_05566_)
  );
  NOR2X1 _12362_ (
    .A(_05542_),
    .B(_05566_),
    .Y(_05463_)
  );
  AOI21X1 _12363_ (
    .A( watchdog_0.wdtcnt_11_ ),
    .B(_05565_),
    .C( watchdog_0.wdtcnt_12_ ),
    .Y(_05567_)
  );
  AND2X1 _12364_ (
    .A(_05491_),
    .B(_05503_),
    .Y(_05568_)
  );
  OR2X1 _12365_ (
    .A(_05567_),
    .B(_05568_),
    .Y(_05569_)
  );
  NOR2X1 _12366_ (
    .A(_05542_),
    .B(_05569_),
    .Y(_05464_)
  );
  OAI21X1 _12367_ (
    .A(_05489_),
    .B(_05490_),
    .C( watchdog_0.wdtcnt_13_ ),
    .Y(_05570_)
  );
  NAND2X1 _12368_ (
    .A(_05491_),
    .B(_05504_),
    .Y(_05571_)
  );
  AOI21X1 _12369_ (
    .A(_05570_),
    .B(_05571_),
    .C(_05542_),
    .Y(_05465_)
  );
  AOI21X1 _12370_ (
    .A( watchdog_0.wdtcnt_13_ ),
    .B(_05568_),
    .C( watchdog_0.wdtcnt_14_ ),
    .Y(_05572_)
  );
  NOR2X1 _12371_ (
    .A(_05492_),
    .B(_05508_),
    .Y(_05573_)
  );
  OR2X1 _12372_ (
    .A(_05572_),
    .B(_05573_),
    .Y(_05574_)
  );
  NOR2X1 _12373_ (
    .A(_05542_),
    .B(_05574_),
    .Y(_05466_)
  );
  XNOR2X1 _12374_ (
    .A( watchdog_0.wdtcnt_15_ ),
    .B(_05573_),
    .Y(_05575_)
  );
  NOR2X1 _12375_ (
    .A(_05542_),
    .B(_05575_),
    .Y(_05467_)
  );
  DFFSR _12376_ (
    .CLK(dco_clk),
    .D(_05443_),
    .Q( clock_module_0.wdt_reset ),
    .R(_05444_),
    .S(1'h1)
  );
  DFFSR _12377_ (
    .CLK(dco_clk),
    .D(_05446_),
    .Q( watchdog_0.wdtctl_0_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12378_ (
    .CLK(dco_clk),
    .D(_05447_),
    .Q( watchdog_0.wdtctl_1_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12379_ (
    .CLK(dco_clk),
    .D(_05448_),
    .Q( watchdog_0.wdtctl_2_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12380_ (
    .CLK(dco_clk),
    .D(_05449_),
    .Q( watchdog_0.wdtctl_4_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12381_ (
    .CLK(dco_clk),
    .D(_05450_),
    .Q( watchdog_0.wdtctl_7_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12382_ (
    .CLK(dco_clk),
    .D(_05451_),
    .Q( sfr_0.ifg1_0_ ),
    .R(_05444_),
    .S(1'h1)
  );
  DFFSR _12383_ (
    .CLK(dco_clk),
    .D(_05452_),
    .Q( watchdog_0.wdtcnt_0_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12384_ (
    .CLK(dco_clk),
    .D(_05453_),
    .Q( watchdog_0.wdtcnt_1_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12385_ (
    .CLK(dco_clk),
    .D(_05454_),
    .Q( watchdog_0.wdtcnt_2_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12386_ (
    .CLK(dco_clk),
    .D(_05455_),
    .Q( watchdog_0.wdtcnt_3_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12387_ (
    .CLK(dco_clk),
    .D(_05456_),
    .Q( watchdog_0.wdtcnt_4_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12388_ (
    .CLK(dco_clk),
    .D(_05457_),
    .Q( watchdog_0.wdtcnt_5_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12389_ (
    .CLK(dco_clk),
    .D(_05458_),
    .Q( watchdog_0.wdtcnt_6_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12390_ (
    .CLK(dco_clk),
    .D(_05459_),
    .Q( watchdog_0.wdtcnt_7_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12391_ (
    .CLK(dco_clk),
    .D(_05460_),
    .Q( watchdog_0.wdtcnt_8_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12392_ (
    .CLK(dco_clk),
    .D(_05461_),
    .Q( watchdog_0.wdtcnt_9_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12393_ (
    .CLK(dco_clk),
    .D(_05462_),
    .Q( watchdog_0.wdtcnt_10_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12394_ (
    .CLK(dco_clk),
    .D(_05463_),
    .Q( watchdog_0.wdtcnt_11_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12395_ (
    .CLK(dco_clk),
    .D(_05464_),
    .Q( watchdog_0.wdtcnt_12_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12396_ (
    .CLK(dco_clk),
    .D(_05465_),
    .Q( watchdog_0.wdtcnt_13_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12397_ (
    .CLK(dco_clk),
    .D(_05466_),
    .Q( watchdog_0.wdtcnt_14_ ),
    .R(_05445_),
    .S(1'h1)
  );
  DFFSR _12398_ (
    .CLK(dco_clk),
    .D(_05467_),
    .Q( watchdog_0.wdtcnt_15_ ),
    .R(_05445_),
    .S(1'h1)
  );
  BUFX2 _12399_ (
    .A(dco_clk),
    .Y(aclk)
  );
  BUFX2 _12400_ (
    .A(_05581_),
    .Y(aclk_en)
  );
  BUFX2 _12401_ (
    .A(_05582_),
    .Y(dbg_freeze)
  );
  BUFX2 _12402_ (
    .A(_05583_),
    .Y(dbg_i2c_sda_out)
  );
  BUFX2 _12403_ (
    .A(1'h1),
    .Y(dbg_uart_txd)
  );
  BUFX2 _12404_ (
    .A(1'h1),
    .Y(dco_enable)
  );
  BUFX2 _12405_ (
    .A(1'h1),
    .Y(dco_wkup)
  );
  BUFX2 _12406_ (
    .A(1'h0),
    .Y(dma_dout_0_)
  );
  BUFX2 _12407_ (
    .A(1'h0),
    .Y(dma_dout_10_)
  );
  BUFX2 _12408_ (
    .A(1'h0),
    .Y(dma_dout_11_)
  );
  BUFX2 _12409_ (
    .A(1'h0),
    .Y(dma_dout_12_)
  );
  BUFX2 _12410_ (
    .A(1'h0),
    .Y(dma_dout_13_)
  );
  BUFX2 _12411_ (
    .A(1'h0),
    .Y(dma_dout_14_)
  );
  BUFX2 _12412_ (
    .A(1'h0),
    .Y(dma_dout_15_)
  );
  BUFX2 _12413_ (
    .A(1'h0),
    .Y(dma_dout_1_)
  );
  BUFX2 _12414_ (
    .A(1'h0),
    .Y(dma_dout_2_)
  );
  BUFX2 _12415_ (
    .A(1'h0),
    .Y(dma_dout_3_)
  );
  BUFX2 _12416_ (
    .A(1'h0),
    .Y(dma_dout_4_)
  );
  BUFX2 _12417_ (
    .A(1'h0),
    .Y(dma_dout_5_)
  );
  BUFX2 _12418_ (
    .A(1'h0),
    .Y(dma_dout_6_)
  );
  BUFX2 _12419_ (
    .A(1'h0),
    .Y(dma_dout_7_)
  );
  BUFX2 _12420_ (
    .A(1'h0),
    .Y(dma_dout_8_)
  );
  BUFX2 _12421_ (
    .A(1'h0),
    .Y(dma_dout_9_)
  );
  BUFX2 _12422_ (
    .A(1'h1),
    .Y(dma_ready)
  );
  BUFX2 _12423_ (
    .A(1'h1),
    .Y(dma_resp)
  );
  BUFX2 _12424_ (
    .A(_05584_),
    .Y(dmem_addr_0_)
  );
  BUFX2 _12425_ (
    .A(_05585_),
    .Y(dmem_addr_10_)
  );
  BUFX2 _12426_ (
    .A(_05586_),
    .Y(dmem_addr_11_)
  );
  BUFX2 _12427_ (
    .A(_05587_),
    .Y(dmem_addr_12_)
  );
  BUFX2 _12428_ (
    .A(_05588_),
    .Y(dmem_addr_1_)
  );
  BUFX2 _12429_ (
    .A(_05589_),
    .Y(dmem_addr_2_)
  );
  BUFX2 _12430_ (
    .A(_05590_),
    .Y(dmem_addr_3_)
  );
  BUFX2 _12431_ (
    .A(_05591_),
    .Y(dmem_addr_4_)
  );
  BUFX2 _12432_ (
    .A(_05592_),
    .Y(dmem_addr_5_)
  );
  BUFX2 _12433_ (
    .A(_05593_),
    .Y(dmem_addr_6_)
  );
  BUFX2 _12434_ (
    .A(_05594_),
    .Y(dmem_addr_7_)
  );
  BUFX2 _12435_ (
    .A(_05595_),
    .Y(dmem_addr_8_)
  );
  BUFX2 _12436_ (
    .A(_05596_),
    .Y(dmem_addr_9_)
  );
  BUFX2 _12437_ (
    .A(_05597_),
    .Y(dmem_cen)
  );
  BUFX2 _12438_ (
    .A(_05598_),
    .Y(dmem_din_0_)
  );
  BUFX2 _12439_ (
    .A(_05599_),
    .Y(dmem_din_10_)
  );
  BUFX2 _12440_ (
    .A(_05600_),
    .Y(dmem_din_11_)
  );
  BUFX2 _12441_ (
    .A(_05601_),
    .Y(dmem_din_12_)
  );
  BUFX2 _12442_ (
    .A(_05602_),
    .Y(dmem_din_13_)
  );
  BUFX2 _12443_ (
    .A(_05603_),
    .Y(dmem_din_14_)
  );
  BUFX2 _12444_ (
    .A(_05604_),
    .Y(dmem_din_15_)
  );
  BUFX2 _12445_ (
    .A(_05605_),
    .Y(dmem_din_1_)
  );
  BUFX2 _12446_ (
    .A(_05606_),
    .Y(dmem_din_2_)
  );
  BUFX2 _12447_ (
    .A(_05607_),
    .Y(dmem_din_3_)
  );
  BUFX2 _12448_ (
    .A(_05608_),
    .Y(dmem_din_4_)
  );
  BUFX2 _12449_ (
    .A(_05609_),
    .Y(dmem_din_5_)
  );
  BUFX2 _12450_ (
    .A(_05610_),
    .Y(dmem_din_6_)
  );
  BUFX2 _12451_ (
    .A(_05611_),
    .Y(dmem_din_7_)
  );
  BUFX2 _12452_ (
    .A(_05612_),
    .Y(dmem_din_8_)
  );
  BUFX2 _12453_ (
    .A(_05613_),
    .Y(dmem_din_9_)
  );
  BUFX2 _12454_ (
    .A(_05614_),
    .Y(dmem_wen_0_)
  );
  BUFX2 _12455_ (
    .A(_05615_),
    .Y(dmem_wen_1_)
  );
  BUFX2 _12456_ (
    .A(_05616_),
    .Y(irq_acc_0_)
  );
  BUFX2 _12457_ (
    .A(_05617_),
    .Y(irq_acc_10_)
  );
  BUFX2 _12458_ (
    .A(_05618_),
    .Y(irq_acc_11_)
  );
  BUFX2 _12459_ (
    .A(_05619_),
    .Y(irq_acc_12_)
  );
  BUFX2 _12460_ (
    .A(_05620_),
    .Y(irq_acc_13_)
  );
  BUFX2 _12461_ (
    .A(_05621_),
    .Y(irq_acc_1_)
  );
  BUFX2 _12462_ (
    .A(_05622_),
    .Y(irq_acc_2_)
  );
  BUFX2 _12463_ (
    .A(_05623_),
    .Y(irq_acc_3_)
  );
  BUFX2 _12464_ (
    .A(_05624_),
    .Y(irq_acc_4_)
  );
  BUFX2 _12465_ (
    .A(_05625_),
    .Y(irq_acc_5_)
  );
  BUFX2 _12466_ (
    .A(_05626_),
    .Y(irq_acc_6_)
  );
  BUFX2 _12467_ (
    .A(_05627_),
    .Y(irq_acc_7_)
  );
  BUFX2 _12468_ (
    .A(_05628_),
    .Y(irq_acc_8_)
  );
  BUFX2 _12469_ (
    .A(_05629_),
    .Y(irq_acc_9_)
  );
  BUFX2 _12470_ (
    .A(1'h1),
    .Y(lfxt_enable)
  );
  BUFX2 _12471_ (
    .A(1'h0),
    .Y(lfxt_wkup)
  );
  BUFX2 _12472_ (
    .A(dco_clk),
    .Y(mclk)
  );
  BUFX2 _12473_ (
    .A(_05630_),
    .Y(per_addr_0_)
  );
  BUFX2 _12474_ (
    .A(_05631_),
    .Y(per_addr_10_)
  );
  BUFX2 _12475_ (
    .A(_05632_),
    .Y(per_addr_11_)
  );
  BUFX2 _12476_ (
    .A(_05633_),
    .Y(per_addr_12_)
  );
  BUFX2 _12477_ (
    .A(1'h0),
    .Y(per_addr_13_)
  );
  BUFX2 _12478_ (
    .A(_05634_),
    .Y(per_addr_1_)
  );
  BUFX2 _12479_ (
    .A(_05635_),
    .Y(per_addr_2_)
  );
  BUFX2 _12480_ (
    .A(_05636_),
    .Y(per_addr_3_)
  );
  BUFX2 _12481_ (
    .A(_05637_),
    .Y(per_addr_4_)
  );
  BUFX2 _12482_ (
    .A(_05638_),
    .Y(per_addr_5_)
  );
  BUFX2 _12483_ (
    .A(_05639_),
    .Y(per_addr_6_)
  );
  BUFX2 _12484_ (
    .A(_05640_),
    .Y(per_addr_7_)
  );
  BUFX2 _12485_ (
    .A(_05641_),
    .Y(per_addr_8_)
  );
  BUFX2 _12486_ (
    .A(_05642_),
    .Y(per_addr_9_)
  );
  BUFX2 _12487_ (
    .A(_05643_),
    .Y(per_din_0_)
  );
  BUFX2 _12488_ (
    .A(_05644_),
    .Y(per_din_10_)
  );
  BUFX2 _12489_ (
    .A(_05645_),
    .Y(per_din_11_)
  );
  BUFX2 _12490_ (
    .A(_05646_),
    .Y(per_din_12_)
  );
  BUFX2 _12491_ (
    .A(_05647_),
    .Y(per_din_13_)
  );
  BUFX2 _12492_ (
    .A(_05648_),
    .Y(per_din_14_)
  );
  BUFX2 _12493_ (
    .A(_05649_),
    .Y(per_din_15_)
  );
  BUFX2 _12494_ (
    .A(_05650_),
    .Y(per_din_1_)
  );
  BUFX2 _12495_ (
    .A(_05651_),
    .Y(per_din_2_)
  );
  BUFX2 _12496_ (
    .A(_05652_),
    .Y(per_din_3_)
  );
  BUFX2 _12497_ (
    .A(_05653_),
    .Y(per_din_4_)
  );
  BUFX2 _12498_ (
    .A(_05654_),
    .Y(per_din_5_)
  );
  BUFX2 _12499_ (
    .A(_05655_),
    .Y(per_din_6_)
  );
  BUFX2 _12500_ (
    .A(_05656_),
    .Y(per_din_7_)
  );
  BUFX2 _12501_ (
    .A(_05657_),
    .Y(per_din_8_)
  );
  BUFX2 _12502_ (
    .A(_05658_),
    .Y(per_din_9_)
  );
  BUFX2 _12503_ (
    .A(_05659_),
    .Y(per_en)
  );
  BUFX2 _12504_ (
    .A(_05660_),
    .Y(per_we_0_)
  );
  BUFX2 _12505_ (
    .A(_05661_),
    .Y(per_we_1_)
  );
  BUFX2 _12506_ (
    .A(_05662_),
    .Y(pmem_addr_0_)
  );
  BUFX2 _12507_ (
    .A(_05663_),
    .Y(pmem_addr_10_)
  );
  BUFX2 _12508_ (
    .A(_05664_),
    .Y(pmem_addr_11_)
  );
  BUFX2 _12509_ (
    .A(_05665_),
    .Y(pmem_addr_12_)
  );
  BUFX2 _12510_ (
    .A(_05666_),
    .Y(pmem_addr_13_)
  );
  BUFX2 _12511_ (
    .A(_05667_),
    .Y(pmem_addr_1_)
  );
  BUFX2 _12512_ (
    .A(_05668_),
    .Y(pmem_addr_2_)
  );
  BUFX2 _12513_ (
    .A(_05669_),
    .Y(pmem_addr_3_)
  );
  BUFX2 _12514_ (
    .A(_05670_),
    .Y(pmem_addr_4_)
  );
  BUFX2 _12515_ (
    .A(_05671_),
    .Y(pmem_addr_5_)
  );
  BUFX2 _12516_ (
    .A(_05672_),
    .Y(pmem_addr_6_)
  );
  BUFX2 _12517_ (
    .A(_05673_),
    .Y(pmem_addr_7_)
  );
  BUFX2 _12518_ (
    .A(_05674_),
    .Y(pmem_addr_8_)
  );
  BUFX2 _12519_ (
    .A(_05675_),
    .Y(pmem_addr_9_)
  );
  BUFX2 _12520_ (
    .A(_05676_),
    .Y(pmem_cen)
  );
  BUFX2 _12521_ (
    .A(_05677_),
    .Y(pmem_din_0_)
  );
  BUFX2 _12522_ (
    .A(_05678_),
    .Y(pmem_din_10_)
  );
  BUFX2 _12523_ (
    .A(_05679_),
    .Y(pmem_din_11_)
  );
  BUFX2 _12524_ (
    .A(_05680_),
    .Y(pmem_din_12_)
  );
  BUFX2 _12525_ (
    .A(_05681_),
    .Y(pmem_din_13_)
  );
  BUFX2 _12526_ (
    .A(_05682_),
    .Y(pmem_din_14_)
  );
  BUFX2 _12527_ (
    .A(_05683_),
    .Y(pmem_din_15_)
  );
  BUFX2 _12528_ (
    .A(_05684_),
    .Y(pmem_din_1_)
  );
  BUFX2 _12529_ (
    .A(_05685_),
    .Y(pmem_din_2_)
  );
  BUFX2 _12530_ (
    .A(_05686_),
    .Y(pmem_din_3_)
  );
  BUFX2 _12531_ (
    .A(_05687_),
    .Y(pmem_din_4_)
  );
  BUFX2 _12532_ (
    .A(_05688_),
    .Y(pmem_din_5_)
  );
  BUFX2 _12533_ (
    .A(_05689_),
    .Y(pmem_din_6_)
  );
  BUFX2 _12534_ (
    .A(_05690_),
    .Y(pmem_din_7_)
  );
  BUFX2 _12535_ (
    .A(_05691_),
    .Y(pmem_din_8_)
  );
  BUFX2 _12536_ (
    .A(_05692_),
    .Y(pmem_din_9_)
  );
  BUFX2 _12537_ (
    .A(_05693_),
    .Y(pmem_wen_0_)
  );
  BUFX2 _12538_ (
    .A(_05694_),
    .Y(pmem_wen_1_)
  );
  BUFX2 _12539_ (
    .A(_05695_),
    .Y(puc_rst)
  );
  BUFX2 _12540_ (
    .A(dco_clk),
    .Y(smclk)
  );
  BUFX2 _12541_ (
    .A(_05696_),
    .Y(smclk_en)
  );
endmodule
